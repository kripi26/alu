magic
tech scmos
timestamp 1701538741
<< polysilicon >>
rect 367 490 384 499
rect 361 452 366 480
rect 393 467 397 468
rect 393 464 405 467
rect 402 452 405 464
rect 361 447 405 452
rect -62 98 -19 105
rect -59 37 -18 44
rect -70 -140 -31 -133
rect -67 -201 -33 -194
rect -70 -393 -34 -386
rect -65 -454 -30 -447
rect -72 -653 -33 -646
rect -58 -714 -28 -707
rect 623 -2036 669 -2032
rect 679 -2063 691 -2059
rect 687 -2078 691 -2063
rect 648 -2084 691 -2078
<< polycontact >>
rect 353 1821 362 1834
rect 472 1753 484 1761
rect 469 1688 482 1700
rect 420 1664 431 1676
rect 394 1639 400 1651
rect 386 1298 395 1303
rect 360 1193 368 1213
rect 440 1188 448 1195
rect 413 1173 425 1180
rect 1165 1166 1172 1171
rect 1185 1120 1191 1124
rect 1227 1072 1235 1079
rect 1203 1043 1207 1056
rect 385 936 390 944
rect 436 796 443 804
rect 404 775 416 782
rect 360 490 367 499
rect 361 480 366 486
rect -71 98 -62 105
rect -68 37 -59 44
rect 577 -112 588 -103
rect -88 -140 -70 -133
rect 591 -163 596 -156
rect -77 -201 -67 -194
rect 660 -307 665 -300
rect 623 -322 630 -314
rect -81 -393 -70 -386
rect -74 -454 -65 -447
rect -80 -653 -72 -646
rect -65 -714 -58 -707
rect 476 -961 493 -951
rect 454 -974 462 -961
rect 527 -991 540 -983
rect 545 -1021 552 -1014
rect 423 -1107 433 -1097
rect 548 -1333 556 -1329
rect 574 -1420 583 -1398
rect 619 -1423 635 -1416
rect 649 -1470 655 -1463
rect 1171 -1535 1177 -1530
rect 1182 -1559 1188 -1552
rect 1227 -1629 1233 -1622
rect 1202 -1676 1209 -1669
rect 548 -1730 557 -1722
rect 588 -1791 597 -1779
rect 643 -1825 649 -1817
rect 616 -2036 623 -2032
rect 641 -2084 648 -2078
<< metal1 >>
rect -449 1899 484 1916
rect 546 1909 555 1970
rect 719 1909 1299 1917
rect -449 -462 -432 1899
rect -389 1821 353 1834
rect -389 -646 -381 1821
rect 472 1761 484 1899
rect -70 1609 -41 1614
rect -28 1609 -22 1674
rect -70 1332 -65 1609
rect 394 1583 400 1639
rect -6 1580 400 1583
rect -2 1551 36 1557
rect -70 1327 -33 1332
rect -70 1010 -65 1327
rect -3 1298 14 1303
rect 28 1275 36 1551
rect 420 1507 431 1664
rect 5 1269 36 1275
rect -70 1005 -32 1010
rect -70 819 -65 1005
rect -1 976 12 981
rect 28 953 36 1269
rect 136 1495 431 1507
rect 136 1068 148 1495
rect 469 1466 482 1688
rect 807 1603 1172 1607
rect 200 1455 482 1466
rect 200 1125 213 1455
rect 334 1298 386 1303
rect 321 1193 360 1213
rect 200 1120 314 1125
rect 314 959 319 1120
rect 413 1068 425 1173
rect 440 1125 448 1188
rect 733 1182 1052 1185
rect 1049 1124 1052 1182
rect 1165 1171 1172 1603
rect 1288 1197 1299 1909
rect 1049 1120 1185 1124
rect 345 976 390 981
rect 7 947 36 953
rect -106 808 -65 819
rect -106 224 -93 808
rect -70 748 -65 808
rect -70 743 -32 748
rect -1 714 9 719
rect 28 691 36 947
rect 385 944 390 976
rect 413 804 425 1056
rect 930 1043 1203 1056
rect 336 796 436 804
rect 930 795 939 1043
rect 694 792 939 795
rect 8 685 15 691
rect 27 685 36 691
rect 404 647 416 775
rect -2 637 416 647
rect -34 490 360 499
rect 1227 491 1235 1072
rect 1461 1063 1498 1066
rect 469 487 1235 491
rect 74 480 361 486
rect 314 291 319 463
rect 329 289 336 448
rect -158 220 702 224
rect -159 211 702 220
rect -159 -52 -143 211
rect -127 -3 -119 185
rect 134 178 142 211
rect -89 98 -71 105
rect 280 92 329 97
rect 336 92 545 97
rect 552 92 588 97
rect -87 37 -68 44
rect -159 -60 58 -52
rect -372 -201 -244 -194
rect -372 -603 -365 -201
rect -195 -612 -187 -140
rect -159 -305 -143 -60
rect 577 -103 588 92
rect 689 -65 702 211
rect -119 -140 -88 -133
rect 280 -146 314 -141
rect 319 -146 527 -141
rect 540 -146 596 -141
rect 591 -156 596 -146
rect -101 -201 -77 -194
rect -159 -313 63 -305
rect -159 -565 -144 -313
rect -99 -393 -81 -386
rect 624 -392 630 -322
rect 282 -399 477 -392
rect 493 -399 630 -392
rect -104 -454 -74 -447
rect 341 -529 351 -399
rect -102 -536 351 -529
rect -159 -573 -82 -565
rect -75 -573 60 -565
rect -389 -653 -80 -646
rect -338 -753 -310 -691
rect -337 -1398 -311 -753
rect -240 -1379 -232 -1363
rect -241 -1538 -232 -1379
rect -195 -1511 -187 -696
rect -175 -713 -163 -653
rect 660 -654 665 -307
rect 930 -313 951 -310
rect 282 -659 665 -654
rect -176 -1093 -163 -713
rect -88 -714 -65 -707
rect 356 -838 370 -753
rect 477 -789 493 -692
rect -29 -846 370 -838
rect 527 -831 540 -691
rect 545 -822 552 -692
rect -29 -847 367 -846
rect -176 -1161 -164 -1093
rect -29 -1142 -21 -847
rect 313 -866 593 -858
rect 790 -866 1356 -858
rect 313 -870 314 -866
rect 302 -979 314 -870
rect 476 -912 477 -898
rect 476 -951 493 -912
rect 395 -974 454 -961
rect 527 -983 540 -915
rect 284 -1107 423 -1097
rect -176 -1166 0 -1161
rect 284 -1162 289 -1107
rect 40 -1165 289 -1162
rect -103 -1194 -29 -1188
rect -21 -1194 7 -1188
rect 527 -1262 540 -991
rect 545 -1014 552 -914
rect 545 -1245 552 -1021
rect 875 -1172 1177 -1168
rect 545 -1253 655 -1245
rect 619 -1262 635 -1261
rect 527 -1274 635 -1262
rect -57 -1304 9 -1299
rect -63 -1480 -57 -1304
rect 36 -1333 548 -1329
rect 114 -1419 574 -1398
rect 619 -1416 635 -1274
rect 649 -1463 655 -1253
rect 649 -1473 655 -1470
rect 643 -1478 655 -1473
rect -57 -1486 7 -1481
rect -195 -1516 -4 -1511
rect 34 -1515 515 -1511
rect 403 -1516 515 -1515
rect -241 -1544 5 -1538
rect -241 -1717 -232 -1544
rect 460 -1610 477 -1609
rect -123 -1623 478 -1610
rect 41 -1694 293 -1691
rect -241 -1723 5 -1717
rect -43 -2105 -36 -1723
rect 282 -2032 293 -1694
rect 460 -1779 477 -1623
rect 507 -1722 515 -1516
rect 507 -1730 548 -1722
rect 460 -1791 588 -1779
rect 643 -1817 649 -1478
rect 892 -1526 1141 -1520
rect 1133 -1552 1141 -1526
rect 1171 -1530 1177 -1172
rect 1345 -1504 1356 -866
rect 1133 -1559 1182 -1552
rect 1202 -1869 1209 -1676
rect 857 -1874 1209 -1869
rect 1227 -2032 1233 -1629
rect 1458 -1638 1485 -1635
rect 282 -2036 616 -2032
rect 755 -2039 1236 -2032
rect 609 -2078 615 -2052
rect 609 -2084 641 -2078
rect 707 -2096 717 -2072
rect 706 -2105 717 -2096
rect -43 -2113 717 -2105
rect 706 -2131 717 -2113
rect 1366 -2131 1373 -1799
rect 706 -2141 1373 -2131
<< m2contact >>
rect 546 1970 555 1985
rect -449 -473 -432 -462
rect -28 1674 -22 1681
rect -50 1579 -45 1584
rect -42 1297 -37 1302
rect 14 1298 19 1303
rect -40 975 -35 980
rect 12 976 17 981
rect 693 1585 700 1596
rect 477 1429 483 1436
rect 329 1298 334 1303
rect 296 1193 321 1213
rect 314 1120 319 1125
rect 136 1056 148 1068
rect 440 1120 448 1125
rect 623 1108 633 1115
rect 413 1056 425 1068
rect 340 976 345 981
rect 314 954 319 959
rect -40 713 -35 718
rect 9 714 14 719
rect 462 968 472 980
rect 329 796 336 804
rect 15 685 27 691
rect 592 725 603 734
rect -13 637 -2 647
rect 373 523 378 529
rect -44 490 -34 499
rect 1364 894 1370 901
rect 66 480 74 486
rect 314 463 319 468
rect 314 286 319 291
rect 329 448 336 457
rect 420 455 426 462
rect 329 280 336 289
rect -127 185 -119 195
rect -98 98 -89 105
rect 329 92 336 97
rect 545 92 552 97
rect -94 37 -87 44
rect -127 -10 -119 -3
rect -195 -140 -187 -131
rect -244 -201 -234 -194
rect -372 -610 -365 -603
rect -127 -140 -119 -133
rect 314 -146 319 -141
rect 527 -146 540 -141
rect -111 -201 -101 -194
rect -110 -393 -99 -386
rect 477 -399 493 -392
rect -109 -454 -104 -447
rect -110 -536 -102 -529
rect -82 -574 -75 -565
rect -195 -619 -187 -612
rect -339 -691 -310 -672
rect -195 -696 -187 -685
rect -240 -1363 -232 -1356
rect -337 -1419 -310 -1398
rect 708 -387 725 -380
rect 477 -692 493 -676
rect -95 -714 -88 -707
rect 356 -753 370 -746
rect 477 -803 493 -789
rect 527 -691 540 -676
rect 545 -692 552 -677
rect 545 -831 552 -822
rect 527 -839 540 -831
rect 302 -870 313 -858
rect 477 -912 493 -898
rect 527 -915 540 -905
rect 380 -974 395 -961
rect 302 -992 314 -979
rect 3 -1136 9 -1131
rect -29 -1150 -21 -1142
rect -111 -1194 -103 -1188
rect -29 -1194 -21 -1188
rect 545 -914 552 -905
rect 740 -1190 753 -1179
rect -63 -1304 -57 -1299
rect -3 -1334 2 -1329
rect 2 -1362 10 -1356
rect 85 -1419 114 -1398
rect 665 -1281 673 -1272
rect -63 -1486 -57 -1480
rect -136 -1623 -123 -1610
rect 4 -1665 10 -1660
rect -3 -1695 2 -1690
rect 805 -1600 818 -1593
rect 655 -1698 667 -1686
rect 773 -1941 784 -1932
rect 659 -2003 665 -1998
rect 609 -2052 615 -2044
rect 707 -2072 717 -2065
<< metal2 >>
rect 294 1970 546 1985
rect -22 1674 283 1681
rect -356 1579 -50 1584
rect -449 -529 -432 -473
rect -372 -1611 -365 -610
rect -356 -707 -349 1579
rect 693 1574 700 1585
rect 623 1565 700 1574
rect 294 1429 477 1436
rect -305 1297 -42 1302
rect 19 1298 329 1303
rect -305 -430 -293 1297
rect -277 1193 296 1212
rect -277 -386 -267 1193
rect 319 1120 440 1125
rect 623 1115 633 1565
rect 623 1099 633 1108
rect 592 1091 633 1099
rect 148 1056 413 1068
rect -244 975 -40 980
rect 17 976 340 981
rect -244 -194 -234 975
rect 437 968 462 980
rect -195 713 -40 718
rect 14 714 74 719
rect -195 45 -188 713
rect -127 637 -13 647
rect -127 195 -119 637
rect -44 202 -34 490
rect 15 419 27 685
rect 66 486 74 714
rect 314 468 319 954
rect 329 457 336 796
rect 592 734 603 1091
rect 592 671 603 725
rect 1364 671 1370 894
rect 592 651 1370 671
rect 592 600 603 651
rect 420 592 603 600
rect 346 523 373 529
rect 420 462 426 592
rect 420 419 426 455
rect 15 412 426 419
rect 15 325 27 412
rect 15 305 424 325
rect -98 196 -34 202
rect -98 105 -89 196
rect -165 98 -98 105
rect -188 37 -94 44
rect -127 -132 -119 -10
rect 120 -16 128 3
rect 120 -22 309 -16
rect -187 -133 -119 -132
rect -187 -140 -127 -133
rect -234 -201 -111 -194
rect 299 -232 309 -22
rect 314 -141 319 286
rect 329 97 336 280
rect 212 -240 309 -232
rect -277 -393 -216 -386
rect -204 -393 -110 -386
rect -339 -447 -293 -430
rect -339 -454 -109 -447
rect -339 -672 -310 -454
rect 299 -488 309 -240
rect 214 -493 309 -488
rect -234 -536 -110 -529
rect -82 -598 -75 -574
rect -195 -685 -187 -619
rect -356 -714 -95 -707
rect -136 -961 -127 -714
rect 299 -746 309 -493
rect 412 -746 424 305
rect 477 -676 493 -399
rect 527 -676 540 -146
rect 545 -677 552 92
rect 708 -746 725 -387
rect 299 -748 356 -746
rect 219 -753 356 -748
rect 370 -752 725 -746
rect 370 -753 724 -752
rect -75 -870 302 -858
rect 477 -898 493 -803
rect 527 -905 540 -839
rect 545 -905 552 -831
rect -136 -974 380 -961
rect -56 -1136 3 -1131
rect -240 -1194 -111 -1188
rect -240 -1356 -232 -1194
rect -63 -1299 -57 -1136
rect -29 -1188 -21 -1150
rect 302 -1272 314 -992
rect 740 -1220 753 -1190
rect 740 -1231 818 -1220
rect 302 -1281 665 -1272
rect -204 -1334 -3 -1329
rect -232 -1362 2 -1356
rect -232 -1363 10 -1362
rect -310 -1419 85 -1398
rect -373 -1623 -136 -1611
rect -63 -1660 -58 -1486
rect -63 -1665 4 -1660
rect 302 -1686 314 -1281
rect 805 -1593 818 -1231
rect 805 -1616 818 -1600
rect 774 -1628 818 -1616
rect -468 -1695 -3 -1690
rect 302 -1698 655 -1686
rect 302 -1707 314 -1698
rect 301 -1998 314 -1707
rect 773 -1932 784 -1628
rect 773 -1956 784 -1941
rect 700 -1971 784 -1956
rect 301 -2003 659 -1998
rect 700 -2015 710 -1971
rect 700 -2025 717 -2015
rect -455 -2052 609 -2044
rect 707 -2065 717 -2025
<< m3contact >>
rect 283 1970 294 1985
rect 283 1674 294 1681
rect -449 -536 -432 -529
rect 283 1429 294 1436
rect 428 968 437 980
rect 341 523 346 529
rect -173 98 -165 105
rect -195 37 -188 45
rect -216 -393 -204 -386
rect -251 -536 -234 -529
rect -82 -608 -75 -598
rect -82 -870 -75 -858
rect -63 -1136 -56 -1131
rect -216 -1334 -204 -1329
rect -478 -1695 -468 -1690
rect -462 -2052 -455 -2044
<< metal3 >>
rect 283 1681 294 1970
rect 283 1436 294 1674
rect 283 980 294 1429
rect 283 968 428 980
rect 283 529 294 968
rect 283 523 341 529
rect -478 98 -173 105
rect -478 -1690 -468 98
rect -462 37 -195 45
rect -462 -2044 -455 37
rect -432 -536 -251 -529
rect -216 -1329 -204 -393
rect -82 -858 -75 -608
rect -82 -1131 -75 -870
rect -82 -1136 -63 -1131
use not  not_7
timestamp 1698771081
transform 1 0 4 0 1 -1695
box -7 -28 41 38
use and  and_1
timestamp 1699973769
transform 1 0 696 0 1 -2034
box -43 -38 74 36
use 3input_AND  3input_AND_1
timestamp 1700474897
transform 1 0 669 0 1 -1775
box -121 -166 219 89
use 4input_AND  4input_AND_2
timestamp 1700476597
transform 1 0 702 0 1 -1396
box -154 -204 219 124
use 4input_OR  4input_OR_1
timestamp 1698909982
transform 1 0 1294 0 1 -1568
box -132 -239 164 71
use 5input_AND  5input_AND_1
timestamp 1700471499
transform 1 0 615 0 1 -921
box -191 -280 263 63
use not  not_6
timestamp 1698771081
transform 1 0 3 0 1 -1516
box -7 -28 41 38
use not  not_5
timestamp 1698771081
transform 1 0 4 0 1 -1334
box -7 -28 41 38
use not  not_4
timestamp 1698771081
transform 1 0 3 0 1 -1166
box -7 -28 41 38
use xnor  xnor_3
timestamp 1700470836
transform 1 0 13 0 1 -733
box -54 -20 299 168
use xnor  xnor_1
timestamp 1700470836
transform 1 0 11 0 1 -220
box -54 -20 299 168
use xnor  xnor_2
timestamp 1700470836
transform 1 0 13 0 1 -473
box -54 -20 299 168
use 4input_AND  4input_AND_0
timestamp 1700476597
transform 1 0 711 0 1 -183
box -154 -204 219 124
use xnor  xnor_0
timestamp 1700470836
transform 1 0 11 0 1 18
box -54 -20 299 168
use and  and_0
timestamp 1699973769
transform 1 0 410 0 1 493
box -43 -38 74 36
use not  not_3
timestamp 1698771081
transform 1 0 -33 0 1 713
box -7 -28 41 38
use 3input_AND  3input_AND_0
timestamp 1700474897
transform 1 0 476 0 1 891
box -121 -166 219 89
use not  not_2
timestamp 1698771081
transform 1 0 -33 0 1 975
box -7 -28 41 38
use 4input_OR  4input_OR_0
timestamp 1698909982
transform 1 0 1297 0 1 1133
box -132 -239 164 71
use not  not_1
timestamp 1698771081
transform 1 0 -35 0 1 1297
box -7 -28 41 38
use 4input_AND  4input_AND_1
timestamp 1700476597
transform 1 0 514 0 1 1312
box -154 -204 219 124
use 5input_AND  5input_AND_0
timestamp 1700471499
transform 1 0 544 0 1 1854
box -191 -280 263 63
use not  not_0
timestamp 1698771081
transform 1 0 -43 0 1 1579
box -7 -28 41 38
<< labels >>
rlabel metal1 -81 100 -81 100 1 a3
rlabel metal1 -80 40 -80 40 1 b3
rlabel metal1 -105 -136 -105 -136 1 a2
rlabel metal1 -88 -197 -88 -197 1 b2
rlabel metal1 -92 -390 -92 -390 1 a1
rlabel metal1 -90 -452 -90 -452 1 b1
rlabel metal1 -89 -650 -89 -650 1 a0
rlabel metal1 -77 -711 -77 -711 1 b0
rlabel metal1 376 215 376 215 1 vdd
rlabel metal2 389 -749 389 -749 1 gnd
rlabel metal1 8 715 9 716 1 b3bar
rlabel m2contact 13 977 14 978 1 b2bar
rlabel m2contact 16 1299 16 1299 1 b1bar
rlabel metal1 4 1581 5 1582 1 b0bar
rlabel metal1 63 -1163 63 -1163 1 a0bar
rlabel metal1 58 -1332 58 -1332 1 a1bar
rlabel metal1 57 -1514 57 -1514 1 a2bar
rlabel metal1 59 -1693 59 -1693 1 a3bar
rlabel metal1 360 95 360 95 1 a3xnorb3
rlabel metal1 369 -143 369 -143 1 a2xnorb2
rlabel metal1 368 -397 368 -397 1 a1xnorb1
rlabel metal1 354 -657 354 -657 1 a0xnorb0
rlabel metal1 816 488 816 488 1 t5
rlabel metal1 935 919 935 919 1 t6
rlabel metal1 956 1183 956 1183 1 t7
rlabel metal1 965 1604 965 1604 1 t8
rlabel metal1 1034 -2035 1034 -2035 1 t1
rlabel metal1 1087 -1873 1087 -1873 1 t2
rlabel metal1 1044 -1525 1044 -1525 1 t3
rlabel metal1 1011 -1170 1011 -1170 1 t4
rlabel metal1 1490 1063 1494 1066 1 out0
rlabel metal1 943 -311 943 -311 1 out1
rlabel metal1 1478 -1638 1482 -1635 1 out2
<< end >>
