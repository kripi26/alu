* SPICE3 file created from alu.ext - technology: scmos
.include TSMC_180nm.txt
.param SUPPLY = 1.8
.param LAMBDA = 0.09u
.param width_P = 8*LAMBDA
.param width_N = 4*LAMBDA
.global gnd vdd

Vdd vdd gnd 1.8
vs0 s0 gnd DC 0
vs1 s1 gnd DC 0
va0 a0 gnd DC 0
va1 a1 gnd DC 0
va2 a2 gnd DC 0
va3 a3 gnd DC 0
vb0 b0 gnd pulse 0 1.8 0ns 100ps 100ps 20ns 40ns
vb1 b1 gnd pulse 0 1.8 0ns 100ps 100ps 20ns 40ns
vb2 b2 gnd pulse 0 1.8 0ns 100ps 100ps 20ns 40ns
vb3 b3 gnd pulse 0 1.8 0ns 100ps 100ps 20ns 40ns


* *and block
* Vdd vdd gnd 1.8
* vs0 s0 gnd DC 1.8
* vs1 s1 gnd DC 1.8
* vb0 b0 gnd DC 1.8
* vb1 b1 gnd DC 1.8
* vb2 b2 gnd DC 1.8
* vb3 b3 gnd DC 1.8
* va0 a0 gnd pulse 0 1.8 0ns 100ps 100ps 20ns 40ns
* va1 a1 gnd pulse 0 1.8 0ns 100ps 100ps 20ns 40ns
* va2 a2 gnd pulse 0 1.8 0ns 100ps 100ps 20ns 40ns
* va3 a3 gnd pulse 0 1.8 0ns 100ps 100ps 20ns 40ns

* * sub block
* Vdd vdd gnd 1.8
* vs0 s0 gnd DC 1.8
* vs1 s1 gnd DC 0
* vb0 a0 gnd DC 1.8
* vb1 a1 gnd DC 1.8
* vb2 a2 gnd DC 1.8
* vb3 a3 gnd DC 1.8
* va0 b0 gnd pulse 0 1.8 0ns 100ps 100ps 20ns 40ns
* va1 b1 gnd pulse 0 1.8 0ns 100ps 100ps 20ns 40ns
* va2 b2 gnd pulse 0 1.8 0ns 100ps 100ps 20ns 40ns
* va3 b3 gnd pulse 0 1.8 0ns 100ps 100ps 20ns 40ns

.option scale=0.09u

M1000 b1out_0 enable_0/and_5/a_n26_14# vdd enable_0/and_5/w_26_9# CMOSP w=7 l=4
+  ad=184 pd=80 as=24003 ps=10478
M1001 vdd b1 enable_0/and_5/a_n26_14# enable_0/and_5/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1002 b1out_0 enable_0/and_5/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=309 pd=102 as=48401 ps=12710
M1003 enable_0/and_5/a_n26_14# enable_0/en vdd enable_0/and_5/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1004 enable_0/and_5/a_n26_n23# enable_0/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1005 enable_0/and_5/a_n26_14# b1 enable_0/and_5/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1006 b3out_0 enable_0/and_7/a_n26_14# vdd enable_0/and_7/w_26_9# CMOSP w=7 l=4
+  ad=184 pd=80 as=0 ps=0
M1007 vdd b3 enable_0/and_7/a_n26_14# enable_0/and_7/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1008 b3out_0 enable_0/and_7/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=309 pd=102 as=0 ps=0
M1009 enable_0/and_7/a_n26_14# enable_0/en vdd enable_0/and_7/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1010 enable_0/and_7/a_n26_n23# enable_0/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1011 enable_0/and_7/a_n26_14# b3 enable_0/and_7/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1012 b2out_0 enable_0/and_6/a_n26_14# vdd enable_0/and_6/w_26_9# CMOSP w=7 l=4
+  ad=184 pd=80 as=0 ps=0
M1013 vdd b2 enable_0/and_6/a_n26_14# enable_0/and_6/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1014 b2out_0 enable_0/and_6/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=309 pd=102 as=0 ps=0
M1015 enable_0/and_6/a_n26_14# enable_0/en vdd enable_0/and_6/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1016 enable_0/and_6/a_n26_n23# enable_0/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1017 enable_0/and_6/a_n26_14# b2 enable_0/and_6/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1018 a0out_0 enable_0/and_0/a_n26_14# vdd enable_0/and_0/w_26_9# CMOSP w=7 l=4
+  ad=184 pd=80 as=0 ps=0
M1019 vdd a0 enable_0/and_0/a_n26_14# enable_0/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1020 a0out_0 enable_0/and_0/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=309 pd=102 as=0 ps=0
M1021 enable_0/and_0/a_n26_14# enable_0/en vdd enable_0/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1022 enable_0/and_0/a_n26_n23# enable_0/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1023 enable_0/and_0/a_n26_14# a0 enable_0/and_0/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1024 a1out_0 enable_0/and_1/a_n26_14# vdd enable_0/and_1/w_26_9# CMOSP w=7 l=4
+  ad=184 pd=80 as=0 ps=0
M1025 vdd a1 enable_0/and_1/a_n26_14# enable_0/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1026 a1out_0 enable_0/and_1/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=309 pd=102 as=0 ps=0
M1027 enable_0/and_1/a_n26_14# enable_0/en vdd enable_0/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1028 enable_0/and_1/a_n26_n23# enable_0/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1029 enable_0/and_1/a_n26_14# a1 enable_0/and_1/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1030 a2out_0 enable_0/and_2/a_n26_14# vdd enable_0/and_2/w_26_9# CMOSP w=7 l=4
+  ad=184 pd=80 as=0 ps=0
M1031 vdd a2 enable_0/and_2/a_n26_14# enable_0/and_2/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1032 a2out_0 enable_0/and_2/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=309 pd=102 as=0 ps=0
M1033 enable_0/and_2/a_n26_14# enable_0/en vdd enable_0/and_2/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1034 enable_0/and_2/a_n26_n23# enable_0/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1035 enable_0/and_2/a_n26_14# a2 enable_0/and_2/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1036 a3out_0 enable_0/and_3/a_n26_14# vdd enable_0/and_3/w_26_9# CMOSP w=7 l=4
+  ad=184 pd=80 as=0 ps=0
M1037 vdd a3 enable_0/and_3/a_n26_14# enable_0/and_3/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1038 a3out_0 enable_0/and_3/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=309 pd=102 as=0 ps=0
M1039 enable_0/and_3/a_n26_14# enable_0/en vdd enable_0/and_3/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1040 enable_0/and_3/a_n26_n23# enable_0/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1041 enable_0/and_3/a_n26_14# a3 enable_0/and_3/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1042 b0out_0 enable_0/and_4/a_n26_14# vdd enable_0/and_4/w_26_9# CMOSP w=7 l=4
+  ad=184 pd=80 as=0 ps=0
M1043 vdd b0 enable_0/and_4/a_n26_14# enable_0/and_4/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1044 b0out_0 enable_0/and_4/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=309 pd=102 as=0 ps=0
M1045 enable_0/and_4/a_n26_14# enable_0/en vdd enable_0/and_4/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1046 enable_0/and_4/a_n26_n23# enable_0/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1047 enable_0/and_4/a_n26_14# b0 enable_0/and_4/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1048 b1out_1 enable_1/and_5/a_n26_14# vdd enable_1/and_5/w_26_9# CMOSP w=7 l=4
+  ad=184 pd=80 as=0 ps=0
M1049 vdd b1 enable_1/and_5/a_n26_14# enable_1/and_5/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1050 b1out_1 enable_1/and_5/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=309 pd=102 as=0 ps=0
M1051 enable_1/and_5/a_n26_14# enable_1/en vdd enable_1/and_5/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1052 enable_1/and_5/a_n26_n23# enable_1/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1053 enable_1/and_5/a_n26_14# b1 enable_1/and_5/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1054 b3out_1 enable_1/and_7/a_n26_14# vdd enable_1/and_7/w_26_9# CMOSP w=7 l=4
+  ad=184 pd=80 as=0 ps=0
M1055 vdd b3 enable_1/and_7/a_n26_14# enable_1/and_7/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1056 b3out_1 enable_1/and_7/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=309 pd=102 as=0 ps=0
M1057 enable_1/and_7/a_n26_14# enable_1/en vdd enable_1/and_7/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1058 enable_1/and_7/a_n26_n23# enable_1/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1059 enable_1/and_7/a_n26_14# b3 enable_1/and_7/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1060 b2out_1 enable_1/and_6/a_n26_14# vdd enable_1/and_6/w_26_9# CMOSP w=7 l=4
+  ad=184 pd=80 as=0 ps=0
M1061 vdd b2 enable_1/and_6/a_n26_14# enable_1/and_6/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1062 b2out_1 enable_1/and_6/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=309 pd=102 as=0 ps=0
M1063 enable_1/and_6/a_n26_14# enable_1/en vdd enable_1/and_6/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1064 enable_1/and_6/a_n26_n23# enable_1/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1065 enable_1/and_6/a_n26_14# b2 enable_1/and_6/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1066 a0_out1 enable_1/and_0/a_n26_14# vdd enable_1/and_0/w_26_9# CMOSP w=7 l=4
+  ad=184 pd=80 as=0 ps=0
M1067 vdd a0 enable_1/and_0/a_n26_14# enable_1/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1068 a0_out1 enable_1/and_0/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=309 pd=102 as=0 ps=0
M1069 enable_1/and_0/a_n26_14# enable_1/en vdd enable_1/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1070 enable_1/and_0/a_n26_n23# enable_1/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1071 enable_1/and_0/a_n26_14# a0 enable_1/and_0/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1072 a1out_1 enable_1/and_1/a_n26_14# vdd enable_1/and_1/w_26_9# CMOSP w=7 l=4
+  ad=184 pd=80 as=0 ps=0
M1073 vdd a1 enable_1/and_1/a_n26_14# enable_1/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1074 a1out_1 enable_1/and_1/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=309 pd=102 as=0 ps=0
M1075 enable_1/and_1/a_n26_14# enable_1/en vdd enable_1/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1076 enable_1/and_1/a_n26_n23# enable_1/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1077 enable_1/and_1/a_n26_14# a1 enable_1/and_1/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1078 a2out_1 enable_1/and_2/a_n26_14# vdd enable_1/and_2/w_26_9# CMOSP w=7 l=4
+  ad=184 pd=80 as=0 ps=0
M1079 vdd a2 enable_1/and_2/a_n26_14# enable_1/and_2/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1080 a2out_1 enable_1/and_2/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=309 pd=102 as=0 ps=0
M1081 enable_1/and_2/a_n26_14# enable_1/en vdd enable_1/and_2/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1082 enable_1/and_2/a_n26_n23# enable_1/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1083 enable_1/and_2/a_n26_14# a2 enable_1/and_2/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1084 a3out_1 enable_1/and_3/a_n26_14# vdd enable_1/and_3/w_26_9# CMOSP w=7 l=4
+  ad=184 pd=80 as=0 ps=0
M1085 vdd a3 enable_1/and_3/a_n26_14# enable_1/and_3/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1086 a3out_1 enable_1/and_3/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=309 pd=102 as=0 ps=0
M1087 enable_1/and_3/a_n26_14# enable_1/en vdd enable_1/and_3/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1088 enable_1/and_3/a_n26_n23# enable_1/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1089 enable_1/and_3/a_n26_14# a3 enable_1/and_3/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1090 b0out_1 enable_1/and_4/a_n26_14# vdd enable_1/and_4/w_26_9# CMOSP w=7 l=4
+  ad=184 pd=80 as=0 ps=0
M1091 vdd b0 enable_1/and_4/a_n26_14# enable_1/and_4/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1092 b0out_1 enable_1/and_4/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=309 pd=102 as=0 ps=0
M1093 enable_1/and_4/a_n26_14# enable_1/en vdd enable_1/and_4/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1094 enable_1/and_4/a_n26_n23# enable_1/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1095 enable_1/and_4/a_n26_14# b0 enable_1/and_4/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1096 b1out_3 enable_3/and_5/a_n26_14# vdd enable_3/and_5/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1097 vdd b1 enable_3/and_5/a_n26_14# enable_3/and_5/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1098 b1out_3 enable_3/and_5/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1099 enable_3/and_5/a_n26_14# enable_3/en vdd enable_3/and_5/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1100 enable_3/and_5/a_n26_n23# enable_3/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1101 enable_3/and_5/a_n26_14# b1 enable_3/and_5/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1102 b3out_3 enable_3/and_7/a_n26_14# vdd enable_3/and_7/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1103 vdd b3 enable_3/and_7/a_n26_14# enable_3/and_7/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1104 b3out_3 enable_3/and_7/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1105 enable_3/and_7/a_n26_14# enable_3/en vdd enable_3/and_7/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1106 enable_3/and_7/a_n26_n23# enable_3/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1107 enable_3/and_7/a_n26_14# b3 enable_3/and_7/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1108 b2out_3 enable_3/and_6/a_n26_14# vdd enable_3/and_6/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1109 vdd b2 enable_3/and_6/a_n26_14# enable_3/and_6/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1110 b2out_3 enable_3/and_6/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1111 enable_3/and_6/a_n26_14# enable_3/en vdd enable_3/and_6/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1112 enable_3/and_6/a_n26_n23# enable_3/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1113 enable_3/and_6/a_n26_14# b2 enable_3/and_6/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1114 a0out_3 enable_3/and_0/a_n26_14# vdd enable_3/and_0/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1115 vdd a0 enable_3/and_0/a_n26_14# enable_3/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1116 a0out_3 enable_3/and_0/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1117 enable_3/and_0/a_n26_14# enable_3/en vdd enable_3/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1118 enable_3/and_0/a_n26_n23# enable_3/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1119 enable_3/and_0/a_n26_14# a0 enable_3/and_0/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1120 a1out_3 enable_3/and_1/a_n26_14# vdd enable_3/and_1/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1121 vdd a1 enable_3/and_1/a_n26_14# enable_3/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1122 a1out_3 enable_3/and_1/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1123 enable_3/and_1/a_n26_14# enable_3/en vdd enable_3/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1124 enable_3/and_1/a_n26_n23# enable_3/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1125 enable_3/and_1/a_n26_14# a1 enable_3/and_1/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1126 a2out_3 enable_3/and_2/a_n26_14# vdd enable_3/and_2/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1127 vdd a2 enable_3/and_2/a_n26_14# enable_3/and_2/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1128 a2out_3 enable_3/and_2/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1129 enable_3/and_2/a_n26_14# enable_3/en vdd enable_3/and_2/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1130 enable_3/and_2/a_n26_n23# enable_3/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1131 enable_3/and_2/a_n26_14# a2 enable_3/and_2/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1132 a3out_3 enable_3/and_3/a_n26_14# vdd enable_3/and_3/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1133 vdd a3 enable_3/and_3/a_n26_14# enable_3/and_3/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1134 a3out_3 enable_3/and_3/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1135 enable_3/and_3/a_n26_14# enable_3/en vdd enable_3/and_3/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1136 enable_3/and_3/a_n26_n23# enable_3/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1137 enable_3/and_3/a_n26_14# a3 enable_3/and_3/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1138 b0out_3 enable_3/and_4/a_n26_14# vdd enable_3/and_4/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1139 vdd b0 enable_3/and_4/a_n26_14# enable_3/and_4/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1140 b0out_3 enable_3/and_4/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1141 enable_3/and_4/a_n26_14# enable_3/en vdd enable_3/and_4/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1142 enable_3/and_4/a_n26_n23# enable_3/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1143 enable_3/and_4/a_n26_14# b0 enable_3/and_4/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1144 b1out_2 enable_2/and_5/a_n26_14# vdd enable_2/and_5/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1145 vdd enable_2/b1 enable_2/and_5/a_n26_14# enable_2/and_5/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1146 b1out_2 enable_2/and_5/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1147 enable_2/and_5/a_n26_14# enable_2/en vdd enable_2/and_5/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1148 enable_2/and_5/a_n26_n23# enable_2/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1149 enable_2/and_5/a_n26_14# enable_2/b1 enable_2/and_5/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1150 b3out_2 enable_2/and_7/a_n26_14# vdd enable_2/and_7/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1151 vdd b3 enable_2/and_7/a_n26_14# enable_2/and_7/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1152 b3out_2 enable_2/and_7/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1153 enable_2/and_7/a_n26_14# enable_2/en vdd enable_2/and_7/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1154 enable_2/and_7/a_n26_n23# enable_2/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1155 enable_2/and_7/a_n26_14# b3 enable_2/and_7/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1156 b2out_2 enable_2/and_6/a_n26_14# vdd enable_2/and_6/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1157 vdd b2 enable_2/and_6/a_n26_14# enable_2/and_6/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1158 b2out_2 enable_2/and_6/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1159 enable_2/and_6/a_n26_14# enable_2/en vdd enable_2/and_6/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1160 enable_2/and_6/a_n26_n23# enable_2/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1161 enable_2/and_6/a_n26_14# b2 enable_2/and_6/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1162 a0out_2 enable_2/and_0/a_n26_14# vdd enable_2/and_0/w_26_9# CMOSP w=7 l=4
+  ad=184 pd=80 as=0 ps=0
M1163 vdd enable_2/a0 enable_2/and_0/a_n26_14# enable_2/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1164 a0out_2 enable_2/and_0/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=309 pd=102 as=0 ps=0
M1165 enable_2/and_0/a_n26_14# enable_2/en vdd enable_2/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1166 enable_2/and_0/a_n26_n23# enable_2/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1167 enable_2/and_0/a_n26_14# enable_2/a0 enable_2/and_0/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1168 a1out_2 enable_2/and_1/a_n26_14# vdd enable_2/and_1/w_26_9# CMOSP w=7 l=4
+  ad=184 pd=80 as=0 ps=0
M1169 vdd a1 enable_2/and_1/a_n26_14# enable_2/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1170 a1out_2 enable_2/and_1/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=309 pd=102 as=0 ps=0
M1171 enable_2/and_1/a_n26_14# enable_2/en vdd enable_2/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1172 enable_2/and_1/a_n26_n23# enable_2/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1173 enable_2/and_1/a_n26_14# a1 enable_2/and_1/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1174 a2out_2 enable_2/and_2/a_n26_14# vdd enable_2/and_2/w_26_9# CMOSP w=7 l=4
+  ad=184 pd=80 as=0 ps=0
M1175 vdd enable_2/a2 enable_2/and_2/a_n26_14# enable_2/and_2/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1176 a2out_2 enable_2/and_2/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=309 pd=102 as=0 ps=0
M1177 enable_2/and_2/a_n26_14# enable_2/en vdd enable_2/and_2/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1178 enable_2/and_2/a_n26_n23# enable_2/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1179 enable_2/and_2/a_n26_14# enable_2/a2 enable_2/and_2/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1180 a3out_2 enable_2/and_3/a_n26_14# vdd enable_2/and_3/w_26_9# CMOSP w=7 l=4
+  ad=184 pd=80 as=0 ps=0
M1181 vdd a3 enable_2/and_3/a_n26_14# enable_2/and_3/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1182 a3out_2 enable_2/and_3/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=309 pd=102 as=0 ps=0
M1183 enable_2/and_3/a_n26_14# enable_2/en vdd enable_2/and_3/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1184 enable_2/and_3/a_n26_n23# enable_2/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1185 enable_2/and_3/a_n26_14# a3 enable_2/and_3/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1186 boout_2 enable_2/and_4/a_n26_14# vdd enable_2/and_4/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1187 vdd b0 enable_2/and_4/a_n26_14# enable_2/and_4/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1188 boout_2 enable_2/and_4/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1189 enable_2/and_4/a_n26_14# enable_2/en vdd enable_2/and_4/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1190 enable_2/and_4/a_n26_n23# enable_2/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1191 enable_2/and_4/a_n26_14# b0 enable_2/and_4/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1192 out0 AND_Block_0/and_0/a_n26_14# vdd AND_Block_0/and_0/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1193 vdd b0out_3 AND_Block_0/and_0/a_n26_14# AND_Block_0/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1194 out0 AND_Block_0/and_0/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1195 AND_Block_0/and_0/a_n26_14# a0out_3 vdd AND_Block_0/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1196 AND_Block_0/and_0/a_n26_n23# a0out_3 gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1197 AND_Block_0/and_0/a_n26_14# b0out_3 AND_Block_0/and_0/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1198 out1 AND_Block_0/and_1/a_n26_14# vdd AND_Block_0/and_1/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1199 vdd b1out_3 AND_Block_0/and_1/a_n26_14# AND_Block_0/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1200 out1 AND_Block_0/and_1/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1201 AND_Block_0/and_1/a_n26_14# a1out_3 vdd AND_Block_0/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1202 AND_Block_0/and_1/a_n26_n23# a1out_3 gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1203 AND_Block_0/and_1/a_n26_14# b1out_3 AND_Block_0/and_1/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1204 out2 AND_Block_0/and_2/a_n26_14# vdd AND_Block_0/and_2/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1205 vdd b2out_3 AND_Block_0/and_2/a_n26_14# AND_Block_0/and_2/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1206 out2 AND_Block_0/and_2/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1207 AND_Block_0/and_2/a_n26_14# a2out_3 vdd AND_Block_0/and_2/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1208 AND_Block_0/and_2/a_n26_n23# a2out_3 gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1209 AND_Block_0/and_2/a_n26_14# b2out_3 AND_Block_0/and_2/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1210 out3 AND_Block_0/and_3/a_n26_14# vdd AND_Block_0/and_3/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1211 vdd b3out_3 AND_Block_0/and_3/a_n26_14# AND_Block_0/and_3/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1212 out3 AND_Block_0/and_3/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1213 AND_Block_0/and_3/a_n26_14# a3out_3 vdd AND_Block_0/and_3/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1214 AND_Block_0/and_3/a_n26_n23# a3out_3 gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1215 AND_Block_0/and_3/a_n26_14# b3out_3 AND_Block_0/and_3/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1216 4bitadder_0/fulladder_0/or_0/a_n15_32# 4bitadder_0/fulladder_0/or_0/a gnd Gnd CMOSN w=16 l=5
+  ad=304 pd=70 as=0 ps=0
M1217 4bitadder_0/c1 4bitadder_0/fulladder_0/or_0/a_n15_32# vdd 4bitadder_0/fulladder_0/or_0/w_58_101# CMOSP w=16 l=6
+  ad=288 pd=68 as=0 ps=0
M1218 gnd 4bitadder_0/fulladder_0/or_0/b 4bitadder_0/fulladder_0/or_0/a_n15_32# Gnd CMOSN w=16 l=5
+  ad=0 pd=0 as=0 ps=0
M1219 4bitadder_0/fulladder_0/or_0/a_n15_32# 4bitadder_0/fulladder_0/or_0/b 4bitadder_0/fulladder_0/or_0/a_n15_107# 4bitadder_0/fulladder_0/or_0/w_n48_101# CMOSP w=16 l=5
+  ad=448 pd=88 as=304 ps=70
M1220 4bitadder_0/c1 4bitadder_0/fulladder_0/or_0/a_n15_32# gnd Gnd CMOSN w=16 l=6
+  ad=320 pd=72 as=0 ps=0
M1221 4bitadder_0/fulladder_0/or_0/a_n15_107# 4bitadder_0/fulladder_0/or_0/a vdd 4bitadder_0/fulladder_0/or_0/w_n48_101# CMOSP w=16 l=5
+  ad=0 pd=0 as=0 ps=0
M1222 4bitadder_0/fulladder_0/or_0/a 4bitadder_0/fulladder_0/and_0/a_n26_14# vdd 4bitadder_0/fulladder_0/and_0/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1223 vdd s0 4bitadder_0/fulladder_0/and_0/a_n26_14# 4bitadder_0/fulladder_0/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1224 4bitadder_0/fulladder_0/or_0/a 4bitadder_0/fulladder_0/and_0/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1225 4bitadder_0/fulladder_0/and_0/a_n26_14# 4bitadder_0/fulladder_0/axorb vdd 4bitadder_0/fulladder_0/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1226 4bitadder_0/fulladder_0/and_0/a_n26_n23# 4bitadder_0/fulladder_0/axorb gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1227 4bitadder_0/fulladder_0/and_0/a_n26_14# s0 4bitadder_0/fulladder_0/and_0/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1228 4bitadder_0/fulladder_0/axorb 4bitadder_0/b0xorM 4bitadder_0/fulladder_0/XOR_0/abar Gnd CMOSN w=11 l=6
+  ad=495 pd=156 as=407 ps=118
M1229 4bitadder_0/fulladder_0/XOR_0/bbar 4bitadder_0/b0xorM gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1230 4bitadder_0/fulladder_0/axorb 4bitadder_0/fulladder_0/XOR_0/bbar 4bitadder_0/fulladder_0/XOR_0/abar 4bitadder_0/fulladder_0/XOR_0/w_62_n20# CMOSP w=12 l=6
+  ad=252 pd=110 as=218 ps=84
M1231 vdd 4bitadder_0/b0xorM 4bitadder_0/fulladder_0/XOR_0/bbar 4bitadder_0/fulladder_0/XOR_0/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1232 4bitadder_0/fulladder_0/axorb 4bitadder_0/b0xorM a0out_0 4bitadder_0/fulladder_0/XOR_0/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1233 4bitadder_0/fulladder_0/XOR_0/abar a0out_0 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1234 vdd a0out_0 4bitadder_0/fulladder_0/XOR_0/abar 4bitadder_0/fulladder_0/XOR_0/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1235 4bitadder_0/fulladder_0/axorb 4bitadder_0/fulladder_0/XOR_0/bbar a0out_0 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1236 4bitadder_0/fulladder_0/or_0/b 4bitadder_0/fulladder_0/and_1/a_n26_14# vdd 4bitadder_0/fulladder_0/and_1/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1237 vdd a0out_0 4bitadder_0/fulladder_0/and_1/a_n26_14# 4bitadder_0/fulladder_0/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1238 4bitadder_0/fulladder_0/or_0/b 4bitadder_0/fulladder_0/and_1/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1239 4bitadder_0/fulladder_0/and_1/a_n26_14# 4bitadder_0/b0xorM vdd 4bitadder_0/fulladder_0/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1240 4bitadder_0/fulladder_0/and_1/a_n26_n23# 4bitadder_0/b0xorM gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1241 4bitadder_0/fulladder_0/and_1/a_n26_14# a0out_0 4bitadder_0/fulladder_0/and_1/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1242 s0_add s0 4bitadder_0/fulladder_0/XOR_1/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1243 4bitadder_0/fulladder_0/XOR_1/bbar s0 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1244 s0_add 4bitadder_0/fulladder_0/XOR_1/bbar 4bitadder_0/fulladder_0/XOR_1/abar 4bitadder_0/fulladder_0/XOR_1/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1245 vdd s0 4bitadder_0/fulladder_0/XOR_1/bbar 4bitadder_0/fulladder_0/XOR_1/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1246 s0_add s0 4bitadder_0/fulladder_0/axorb 4bitadder_0/fulladder_0/XOR_1/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1247 4bitadder_0/fulladder_0/XOR_1/abar 4bitadder_0/fulladder_0/axorb gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1248 vdd 4bitadder_0/fulladder_0/axorb 4bitadder_0/fulladder_0/XOR_1/abar 4bitadder_0/fulladder_0/XOR_1/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1249 s0_add 4bitadder_0/fulladder_0/XOR_1/bbar 4bitadder_0/fulladder_0/axorb Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1250 4bitadder_0/fulladder_1/or_0/a_n15_32# 4bitadder_0/fulladder_1/or_0/a gnd Gnd CMOSN w=16 l=5
+  ad=304 pd=70 as=0 ps=0
M1251 4bitadder_0/c2 4bitadder_0/fulladder_1/or_0/a_n15_32# vdd 4bitadder_0/fulladder_1/or_0/w_58_101# CMOSP w=16 l=6
+  ad=288 pd=68 as=0 ps=0
M1252 gnd 4bitadder_0/fulladder_1/or_0/b 4bitadder_0/fulladder_1/or_0/a_n15_32# Gnd CMOSN w=16 l=5
+  ad=0 pd=0 as=0 ps=0
M1253 4bitadder_0/fulladder_1/or_0/a_n15_32# 4bitadder_0/fulladder_1/or_0/b 4bitadder_0/fulladder_1/or_0/a_n15_107# 4bitadder_0/fulladder_1/or_0/w_n48_101# CMOSP w=16 l=5
+  ad=448 pd=88 as=304 ps=70
M1254 4bitadder_0/c2 4bitadder_0/fulladder_1/or_0/a_n15_32# gnd Gnd CMOSN w=16 l=6
+  ad=320 pd=72 as=0 ps=0
M1255 4bitadder_0/fulladder_1/or_0/a_n15_107# 4bitadder_0/fulladder_1/or_0/a vdd 4bitadder_0/fulladder_1/or_0/w_n48_101# CMOSP w=16 l=5
+  ad=0 pd=0 as=0 ps=0
M1256 4bitadder_0/fulladder_1/or_0/a 4bitadder_0/fulladder_1/and_0/a_n26_14# vdd 4bitadder_0/fulladder_1/and_0/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1257 vdd 4bitadder_0/c1 4bitadder_0/fulladder_1/and_0/a_n26_14# 4bitadder_0/fulladder_1/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1258 4bitadder_0/fulladder_1/or_0/a 4bitadder_0/fulladder_1/and_0/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1259 4bitadder_0/fulladder_1/and_0/a_n26_14# 4bitadder_0/fulladder_1/axorb vdd 4bitadder_0/fulladder_1/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1260 4bitadder_0/fulladder_1/and_0/a_n26_n23# 4bitadder_0/fulladder_1/axorb gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1261 4bitadder_0/fulladder_1/and_0/a_n26_14# 4bitadder_0/c1 4bitadder_0/fulladder_1/and_0/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1262 4bitadder_0/fulladder_1/axorb 4bitadder_0/XOR_1/out 4bitadder_0/fulladder_1/XOR_0/abar Gnd CMOSN w=11 l=6
+  ad=495 pd=156 as=407 ps=118
M1263 4bitadder_0/fulladder_1/XOR_0/bbar 4bitadder_0/XOR_1/out gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1264 4bitadder_0/fulladder_1/axorb 4bitadder_0/fulladder_1/XOR_0/bbar 4bitadder_0/fulladder_1/XOR_0/abar 4bitadder_0/fulladder_1/XOR_0/w_62_n20# CMOSP w=12 l=6
+  ad=252 pd=110 as=218 ps=84
M1265 vdd 4bitadder_0/XOR_1/out 4bitadder_0/fulladder_1/XOR_0/bbar 4bitadder_0/fulladder_1/XOR_0/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1266 4bitadder_0/fulladder_1/axorb 4bitadder_0/XOR_1/out a1out_0 4bitadder_0/fulladder_1/XOR_0/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1267 4bitadder_0/fulladder_1/XOR_0/abar a1out_0 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1268 vdd a1out_0 4bitadder_0/fulladder_1/XOR_0/abar 4bitadder_0/fulladder_1/XOR_0/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1269 4bitadder_0/fulladder_1/axorb 4bitadder_0/fulladder_1/XOR_0/bbar a1out_0 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1270 4bitadder_0/fulladder_1/or_0/b 4bitadder_0/fulladder_1/and_1/a_n26_14# vdd 4bitadder_0/fulladder_1/and_1/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1271 vdd a1out_0 4bitadder_0/fulladder_1/and_1/a_n26_14# 4bitadder_0/fulladder_1/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1272 4bitadder_0/fulladder_1/or_0/b 4bitadder_0/fulladder_1/and_1/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1273 4bitadder_0/fulladder_1/and_1/a_n26_14# 4bitadder_0/XOR_1/out vdd 4bitadder_0/fulladder_1/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1274 4bitadder_0/fulladder_1/and_1/a_n26_n23# 4bitadder_0/XOR_1/out gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1275 4bitadder_0/fulladder_1/and_1/a_n26_14# a1out_0 4bitadder_0/fulladder_1/and_1/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1276 s1_add 4bitadder_0/c1 4bitadder_0/fulladder_1/XOR_1/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1277 4bitadder_0/fulladder_1/XOR_1/bbar 4bitadder_0/c1 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1278 s1_add 4bitadder_0/fulladder_1/XOR_1/bbar 4bitadder_0/fulladder_1/XOR_1/abar 4bitadder_0/fulladder_1/XOR_1/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1279 vdd 4bitadder_0/c1 4bitadder_0/fulladder_1/XOR_1/bbar 4bitadder_0/fulladder_1/XOR_1/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1280 s1_add 4bitadder_0/c1 4bitadder_0/fulladder_1/axorb 4bitadder_0/fulladder_1/XOR_1/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1281 4bitadder_0/fulladder_1/XOR_1/abar 4bitadder_0/fulladder_1/axorb gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1282 vdd 4bitadder_0/fulladder_1/axorb 4bitadder_0/fulladder_1/XOR_1/abar 4bitadder_0/fulladder_1/XOR_1/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1283 s1_add 4bitadder_0/fulladder_1/XOR_1/bbar 4bitadder_0/fulladder_1/axorb Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1284 4bitadder_0/fulladder_2/or_0/a_n15_32# 4bitadder_0/fulladder_2/or_0/a gnd Gnd CMOSN w=16 l=5
+  ad=304 pd=70 as=0 ps=0
M1285 4bitadder_0/c3 4bitadder_0/fulladder_2/or_0/a_n15_32# vdd 4bitadder_0/fulladder_2/or_0/w_58_101# CMOSP w=16 l=6
+  ad=288 pd=68 as=0 ps=0
M1286 gnd 4bitadder_0/fulladder_2/or_0/b 4bitadder_0/fulladder_2/or_0/a_n15_32# Gnd CMOSN w=16 l=5
+  ad=0 pd=0 as=0 ps=0
M1287 4bitadder_0/fulladder_2/or_0/a_n15_32# 4bitadder_0/fulladder_2/or_0/b 4bitadder_0/fulladder_2/or_0/a_n15_107# 4bitadder_0/fulladder_2/or_0/w_n48_101# CMOSP w=16 l=5
+  ad=448 pd=88 as=304 ps=70
M1288 4bitadder_0/c3 4bitadder_0/fulladder_2/or_0/a_n15_32# gnd Gnd CMOSN w=16 l=6
+  ad=320 pd=72 as=0 ps=0
M1289 4bitadder_0/fulladder_2/or_0/a_n15_107# 4bitadder_0/fulladder_2/or_0/a vdd 4bitadder_0/fulladder_2/or_0/w_n48_101# CMOSP w=16 l=5
+  ad=0 pd=0 as=0 ps=0
M1290 4bitadder_0/fulladder_2/or_0/a 4bitadder_0/fulladder_2/and_0/a_n26_14# vdd 4bitadder_0/fulladder_2/and_0/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1291 vdd 4bitadder_0/c2 4bitadder_0/fulladder_2/and_0/a_n26_14# 4bitadder_0/fulladder_2/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1292 4bitadder_0/fulladder_2/or_0/a 4bitadder_0/fulladder_2/and_0/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1293 4bitadder_0/fulladder_2/and_0/a_n26_14# 4bitadder_0/fulladder_2/axorb vdd 4bitadder_0/fulladder_2/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1294 4bitadder_0/fulladder_2/and_0/a_n26_n23# 4bitadder_0/fulladder_2/axorb gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1295 4bitadder_0/fulladder_2/and_0/a_n26_14# 4bitadder_0/c2 4bitadder_0/fulladder_2/and_0/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1296 4bitadder_0/fulladder_2/axorb 4bitadder_0/XOR_2/out 4bitadder_0/fulladder_2/XOR_0/abar Gnd CMOSN w=11 l=6
+  ad=495 pd=156 as=407 ps=118
M1297 4bitadder_0/fulladder_2/XOR_0/bbar 4bitadder_0/XOR_2/out gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1298 4bitadder_0/fulladder_2/axorb 4bitadder_0/fulladder_2/XOR_0/bbar 4bitadder_0/fulladder_2/XOR_0/abar 4bitadder_0/fulladder_2/XOR_0/w_62_n20# CMOSP w=12 l=6
+  ad=252 pd=110 as=218 ps=84
M1299 vdd 4bitadder_0/XOR_2/out 4bitadder_0/fulladder_2/XOR_0/bbar 4bitadder_0/fulladder_2/XOR_0/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1300 4bitadder_0/fulladder_2/axorb 4bitadder_0/XOR_2/out a2out_0 4bitadder_0/fulladder_2/XOR_0/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1301 4bitadder_0/fulladder_2/XOR_0/abar a2out_0 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1302 vdd a2out_0 4bitadder_0/fulladder_2/XOR_0/abar 4bitadder_0/fulladder_2/XOR_0/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1303 4bitadder_0/fulladder_2/axorb 4bitadder_0/fulladder_2/XOR_0/bbar a2out_0 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1304 4bitadder_0/fulladder_2/or_0/b 4bitadder_0/fulladder_2/and_1/a_n26_14# vdd 4bitadder_0/fulladder_2/and_1/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1305 vdd a2out_0 4bitadder_0/fulladder_2/and_1/a_n26_14# 4bitadder_0/fulladder_2/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1306 4bitadder_0/fulladder_2/or_0/b 4bitadder_0/fulladder_2/and_1/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1307 4bitadder_0/fulladder_2/and_1/a_n26_14# 4bitadder_0/XOR_2/out vdd 4bitadder_0/fulladder_2/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1308 4bitadder_0/fulladder_2/and_1/a_n26_n23# 4bitadder_0/XOR_2/out gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1309 4bitadder_0/fulladder_2/and_1/a_n26_14# a2out_0 4bitadder_0/fulladder_2/and_1/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1310 s2_add 4bitadder_0/c2 4bitadder_0/fulladder_2/XOR_1/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1311 4bitadder_0/fulladder_2/XOR_1/bbar 4bitadder_0/c2 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1312 s2_add 4bitadder_0/fulladder_2/XOR_1/bbar 4bitadder_0/fulladder_2/XOR_1/abar 4bitadder_0/fulladder_2/XOR_1/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1313 vdd 4bitadder_0/c2 4bitadder_0/fulladder_2/XOR_1/bbar 4bitadder_0/fulladder_2/XOR_1/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1314 s2_add 4bitadder_0/c2 4bitadder_0/fulladder_2/axorb 4bitadder_0/fulladder_2/XOR_1/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1315 4bitadder_0/fulladder_2/XOR_1/abar 4bitadder_0/fulladder_2/axorb gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1316 vdd 4bitadder_0/fulladder_2/axorb 4bitadder_0/fulladder_2/XOR_1/abar 4bitadder_0/fulladder_2/XOR_1/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1317 s2_add 4bitadder_0/fulladder_2/XOR_1/bbar 4bitadder_0/fulladder_2/axorb Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1318 4bitadder_0/fulladder_3/or_0/a_n15_32# 4bitadder_0/fulladder_3/or_0/a gnd Gnd CMOSN w=16 l=5
+  ad=304 pd=70 as=0 ps=0
M1319 fc_add 4bitadder_0/fulladder_3/or_0/a_n15_32# vdd 4bitadder_0/fulladder_3/or_0/w_58_101# CMOSP w=16 l=6
+  ad=288 pd=68 as=0 ps=0
M1320 gnd 4bitadder_0/fulladder_3/or_0/b 4bitadder_0/fulladder_3/or_0/a_n15_32# Gnd CMOSN w=16 l=5
+  ad=0 pd=0 as=0 ps=0
M1321 4bitadder_0/fulladder_3/or_0/a_n15_32# 4bitadder_0/fulladder_3/or_0/b 4bitadder_0/fulladder_3/or_0/a_n15_107# 4bitadder_0/fulladder_3/or_0/w_n48_101# CMOSP w=16 l=5
+  ad=448 pd=88 as=304 ps=70
M1322 fc_add 4bitadder_0/fulladder_3/or_0/a_n15_32# gnd Gnd CMOSN w=16 l=6
+  ad=320 pd=72 as=0 ps=0
M1323 4bitadder_0/fulladder_3/or_0/a_n15_107# 4bitadder_0/fulladder_3/or_0/a vdd 4bitadder_0/fulladder_3/or_0/w_n48_101# CMOSP w=16 l=5
+  ad=0 pd=0 as=0 ps=0
M1324 4bitadder_0/fulladder_3/or_0/a 4bitadder_0/fulladder_3/and_0/a_n26_14# vdd 4bitadder_0/fulladder_3/and_0/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1325 vdd 4bitadder_0/c3 4bitadder_0/fulladder_3/and_0/a_n26_14# 4bitadder_0/fulladder_3/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1326 4bitadder_0/fulladder_3/or_0/a 4bitadder_0/fulladder_3/and_0/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1327 4bitadder_0/fulladder_3/and_0/a_n26_14# 4bitadder_0/fulladder_3/axorb vdd 4bitadder_0/fulladder_3/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1328 4bitadder_0/fulladder_3/and_0/a_n26_n23# 4bitadder_0/fulladder_3/axorb gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1329 4bitadder_0/fulladder_3/and_0/a_n26_14# 4bitadder_0/c3 4bitadder_0/fulladder_3/and_0/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1330 4bitadder_0/fulladder_3/axorb 4bitadder_0/XOR_3/out 4bitadder_0/fulladder_3/XOR_0/abar Gnd CMOSN w=11 l=6
+  ad=495 pd=156 as=407 ps=118
M1331 4bitadder_0/fulladder_3/XOR_0/bbar 4bitadder_0/XOR_3/out gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1332 4bitadder_0/fulladder_3/axorb 4bitadder_0/fulladder_3/XOR_0/bbar 4bitadder_0/fulladder_3/XOR_0/abar 4bitadder_0/fulladder_3/XOR_0/w_62_n20# CMOSP w=12 l=6
+  ad=252 pd=110 as=218 ps=84
M1333 vdd 4bitadder_0/XOR_3/out 4bitadder_0/fulladder_3/XOR_0/bbar 4bitadder_0/fulladder_3/XOR_0/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1334 4bitadder_0/fulladder_3/axorb 4bitadder_0/XOR_3/out a3out_0 4bitadder_0/fulladder_3/XOR_0/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1335 4bitadder_0/fulladder_3/XOR_0/abar a3out_0 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1336 vdd a3out_0 4bitadder_0/fulladder_3/XOR_0/abar 4bitadder_0/fulladder_3/XOR_0/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1337 4bitadder_0/fulladder_3/axorb 4bitadder_0/fulladder_3/XOR_0/bbar a3out_0 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1338 4bitadder_0/fulladder_3/or_0/b 4bitadder_0/fulladder_3/and_1/a_n26_14# vdd 4bitadder_0/fulladder_3/and_1/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1339 vdd a3out_0 4bitadder_0/fulladder_3/and_1/a_n26_14# 4bitadder_0/fulladder_3/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1340 4bitadder_0/fulladder_3/or_0/b 4bitadder_0/fulladder_3/and_1/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1341 4bitadder_0/fulladder_3/and_1/a_n26_14# 4bitadder_0/XOR_3/out vdd 4bitadder_0/fulladder_3/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1342 4bitadder_0/fulladder_3/and_1/a_n26_n23# 4bitadder_0/XOR_3/out gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1343 4bitadder_0/fulladder_3/and_1/a_n26_14# a3out_0 4bitadder_0/fulladder_3/and_1/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1344 s3_add 4bitadder_0/c3 4bitadder_0/fulladder_3/XOR_1/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1345 4bitadder_0/fulladder_3/XOR_1/bbar 4bitadder_0/c3 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1346 s3_add 4bitadder_0/fulladder_3/XOR_1/bbar 4bitadder_0/fulladder_3/XOR_1/abar 4bitadder_0/fulladder_3/XOR_1/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1347 vdd 4bitadder_0/c3 4bitadder_0/fulladder_3/XOR_1/bbar 4bitadder_0/fulladder_3/XOR_1/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1348 s3_add 4bitadder_0/c3 4bitadder_0/fulladder_3/axorb 4bitadder_0/fulladder_3/XOR_1/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1349 4bitadder_0/fulladder_3/XOR_1/abar 4bitadder_0/fulladder_3/axorb gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1350 vdd 4bitadder_0/fulladder_3/axorb 4bitadder_0/fulladder_3/XOR_1/abar 4bitadder_0/fulladder_3/XOR_1/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1351 s3_add 4bitadder_0/fulladder_3/XOR_1/bbar 4bitadder_0/fulladder_3/axorb Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1352 4bitadder_0/b0xorM s0 4bitadder_0/XOR_0/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1353 4bitadder_0/XOR_0/bbar s0 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1354 4bitadder_0/b0xorM 4bitadder_0/XOR_0/bbar 4bitadder_0/XOR_0/abar 4bitadder_0/XOR_0/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1355 vdd s0 4bitadder_0/XOR_0/bbar 4bitadder_0/XOR_0/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1356 4bitadder_0/b0xorM s0 b0out_0 4bitadder_0/XOR_0/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1357 4bitadder_0/XOR_0/abar b0out_0 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1358 vdd b0out_0 4bitadder_0/XOR_0/abar 4bitadder_0/XOR_0/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1359 4bitadder_0/b0xorM 4bitadder_0/XOR_0/bbar b0out_0 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1360 4bitadder_0/XOR_1/out s0 4bitadder_0/XOR_1/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1361 4bitadder_0/XOR_1/bbar s0 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1362 4bitadder_0/XOR_1/out 4bitadder_0/XOR_1/bbar 4bitadder_0/XOR_1/abar 4bitadder_0/XOR_1/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1363 vdd s0 4bitadder_0/XOR_1/bbar 4bitadder_0/XOR_1/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1364 4bitadder_0/XOR_1/out s0 b1out_0 4bitadder_0/XOR_1/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1365 4bitadder_0/XOR_1/abar b1out_0 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1366 vdd b1out_0 4bitadder_0/XOR_1/abar 4bitadder_0/XOR_1/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1367 4bitadder_0/XOR_1/out 4bitadder_0/XOR_1/bbar b1out_0 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1368 4bitadder_0/XOR_2/out s0 4bitadder_0/XOR_2/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1369 4bitadder_0/XOR_2/bbar s0 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1370 4bitadder_0/XOR_2/out 4bitadder_0/XOR_2/bbar 4bitadder_0/XOR_2/abar 4bitadder_0/XOR_2/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1371 vdd s0 4bitadder_0/XOR_2/bbar 4bitadder_0/XOR_2/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1372 4bitadder_0/XOR_2/out s0 b2out_0 4bitadder_0/XOR_2/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1373 4bitadder_0/XOR_2/abar b2out_0 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1374 vdd b2out_0 4bitadder_0/XOR_2/abar 4bitadder_0/XOR_2/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1375 4bitadder_0/XOR_2/out 4bitadder_0/XOR_2/bbar b2out_0 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1376 4bitadder_0/XOR_3/out s0 4bitadder_0/XOR_3/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1377 4bitadder_0/XOR_3/bbar s0 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1378 4bitadder_0/XOR_3/out 4bitadder_0/XOR_3/bbar 4bitadder_0/XOR_3/abar 4bitadder_0/XOR_3/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1379 vdd s0 4bitadder_0/XOR_3/bbar 4bitadder_0/XOR_3/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1380 4bitadder_0/XOR_3/out s0 b3out_0 4bitadder_0/XOR_3/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1381 4bitadder_0/XOR_3/abar b3out_0 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1382 vdd b3out_0 4bitadder_0/XOR_3/abar 4bitadder_0/XOR_3/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1383 4bitadder_0/XOR_3/out 4bitadder_0/XOR_3/bbar b3out_0 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1384 comparator_0/b0bar boout_2 vdd comparator_0/not_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1385 comparator_0/b0bar boout_2 gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1386 comparator_0/b1bar b1out_2 vdd comparator_0/not_1/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1387 comparator_0/b1bar b1out_2 gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1388 agb comparator_0/4input_OR_0/y vdd comparator_0/4input_OR_0/NOT_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1389 agb comparator_0/4input_OR_0/y gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1390 vdd comparator_0/t8 comparator_0/4input_OR_0/a_n52_24# comparator_0/4input_OR_0/w_n58_n43# CMOSP w=14 l=5
+  ad=0 pd=0 as=126 ps=46
M1391 comparator_0/4input_OR_0/y comparator_0/t8 gnd Gnd CMOSN w=16 l=7
+  ad=704 pd=216 as=0 ps=0
M1392 comparator_0/4input_OR_0/a_n52_4# comparator_0/t6 comparator_0/4input_OR_0/a_n52_n15# comparator_0/4input_OR_0/w_n58_n43# CMOSP w=14 l=5
+  ad=210 pd=58 as=196 ps=56
M1393 comparator_0/4input_OR_0/y comparator_0/t5 gnd Gnd CMOSN w=16 l=7
+  ad=0 pd=0 as=0 ps=0
M1394 comparator_0/4input_OR_0/y comparator_0/t7 gnd Gnd CMOSN w=16 l=7
+  ad=0 pd=0 as=0 ps=0
M1395 comparator_0/4input_OR_0/a_n52_24# comparator_0/t7 comparator_0/4input_OR_0/a_n52_4# comparator_0/4input_OR_0/w_n58_n43# CMOSP w=14 l=5
+  ad=0 pd=0 as=0 ps=0
M1396 comparator_0/4input_OR_0/a_n52_n15# comparator_0/t5 comparator_0/4input_OR_0/y comparator_0/4input_OR_0/w_n58_n43# CMOSP w=14 l=5
+  ad=0 pd=0 as=238 ps=62
M1397 comparator_0/4input_OR_0/y comparator_0/t6 gnd Gnd CMOSN w=16 l=7
+  ad=0 pd=0 as=0 ps=0
M1398 comparator_0/b2bar b2out_2 vdd comparator_0/not_2/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1399 comparator_0/b2bar b2out_2 gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1400 comparator_0/a3xnorb3 comparator_0/xnor_0/not_0/in vdd comparator_0/xnor_0/not_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1401 comparator_0/a3xnorb3 comparator_0/xnor_0/not_0/in gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1402 comparator_0/xnor_0/not_0/in comparator_0/b3 comparator_0/xnor_0/XOR_0/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1403 comparator_0/xnor_0/XOR_0/bbar comparator_0/b3 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1404 comparator_0/xnor_0/not_0/in comparator_0/xnor_0/XOR_0/bbar comparator_0/xnor_0/XOR_0/abar comparator_0/xnor_0/XOR_0/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1405 vdd comparator_0/b3 comparator_0/xnor_0/XOR_0/bbar comparator_0/xnor_0/XOR_0/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1406 comparator_0/xnor_0/not_0/in comparator_0/b3 a3out_2 comparator_0/xnor_0/XOR_0/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1407 comparator_0/xnor_0/XOR_0/abar a3out_2 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1408 vdd a3out_2 comparator_0/xnor_0/XOR_0/abar comparator_0/xnor_0/XOR_0/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1409 comparator_0/xnor_0/not_0/in comparator_0/xnor_0/XOR_0/bbar a3out_2 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1410 comparator_0/b3bar comparator_0/b3 vdd comparator_0/not_3/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1411 comparator_0/b3bar comparator_0/b3 gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1412 comparator_0/a2xnorb2 comparator_0/xnor_1/not_0/in vdd comparator_0/xnor_1/not_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1413 comparator_0/a2xnorb2 comparator_0/xnor_1/not_0/in gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1414 comparator_0/xnor_1/not_0/in b2out_2 comparator_0/xnor_1/XOR_0/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1415 comparator_0/xnor_1/XOR_0/bbar b2out_2 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1416 comparator_0/xnor_1/not_0/in comparator_0/xnor_1/XOR_0/bbar comparator_0/xnor_1/XOR_0/abar comparator_0/xnor_1/XOR_0/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1417 vdd b2out_2 comparator_0/xnor_1/XOR_0/bbar comparator_0/xnor_1/XOR_0/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1418 comparator_0/xnor_1/not_0/in b2out_2 a2out_2 comparator_0/xnor_1/XOR_0/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1419 comparator_0/xnor_1/XOR_0/abar a2out_2 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1420 vdd a2out_2 comparator_0/xnor_1/XOR_0/abar comparator_0/xnor_1/XOR_0/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1421 comparator_0/xnor_1/not_0/in comparator_0/xnor_1/XOR_0/bbar a2out_2 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1422 comparator_0/a0bar a0out_2 vdd comparator_0/not_4/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1423 comparator_0/a0bar a0out_2 gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1424 bga comparator_0/4input_OR_1/y vdd comparator_0/4input_OR_1/NOT_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1425 bga comparator_0/4input_OR_1/y gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1426 vdd comparator_0/t4 comparator_0/4input_OR_1/a_n52_24# comparator_0/4input_OR_1/w_n58_n43# CMOSP w=14 l=5
+  ad=0 pd=0 as=126 ps=46
M1427 comparator_0/4input_OR_1/y comparator_0/t4 gnd Gnd CMOSN w=16 l=7
+  ad=704 pd=216 as=0 ps=0
M1428 comparator_0/4input_OR_1/a_n52_4# comparator_0/t2 comparator_0/4input_OR_1/a_n52_n15# comparator_0/4input_OR_1/w_n58_n43# CMOSP w=14 l=5
+  ad=210 pd=58 as=196 ps=56
M1429 comparator_0/4input_OR_1/y comparator_0/t1 gnd Gnd CMOSN w=16 l=7
+  ad=0 pd=0 as=0 ps=0
M1430 comparator_0/4input_OR_1/y comparator_0/t3 gnd Gnd CMOSN w=16 l=7
+  ad=0 pd=0 as=0 ps=0
M1431 comparator_0/4input_OR_1/a_n52_24# comparator_0/t3 comparator_0/4input_OR_1/a_n52_4# comparator_0/4input_OR_1/w_n58_n43# CMOSP w=14 l=5
+  ad=0 pd=0 as=0 ps=0
M1432 comparator_0/4input_OR_1/a_n52_n15# comparator_0/t1 comparator_0/4input_OR_1/y comparator_0/4input_OR_1/w_n58_n43# CMOSP w=14 l=5
+  ad=0 pd=0 as=238 ps=62
M1433 comparator_0/4input_OR_1/y comparator_0/t2 gnd Gnd CMOSN w=16 l=7
+  ad=0 pd=0 as=0 ps=0
M1434 comparator_0/a1xnorb1 comparator_0/xnor_2/not_0/in vdd comparator_0/xnor_2/not_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1435 comparator_0/a1xnorb1 comparator_0/xnor_2/not_0/in gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1436 comparator_0/xnor_2/not_0/in b1out_2 comparator_0/xnor_2/XOR_0/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1437 comparator_0/xnor_2/XOR_0/bbar b1out_2 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1438 comparator_0/xnor_2/not_0/in comparator_0/xnor_2/XOR_0/bbar comparator_0/xnor_2/XOR_0/abar comparator_0/xnor_2/XOR_0/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1439 vdd b1out_2 comparator_0/xnor_2/XOR_0/bbar comparator_0/xnor_2/XOR_0/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1440 comparator_0/xnor_2/not_0/in b1out_2 a1out_2 comparator_0/xnor_2/XOR_0/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1441 comparator_0/xnor_2/XOR_0/abar a1out_2 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1442 vdd a1out_2 comparator_0/xnor_2/XOR_0/abar comparator_0/xnor_2/XOR_0/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1443 comparator_0/xnor_2/not_0/in comparator_0/xnor_2/XOR_0/bbar a1out_2 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1444 comparator_0/a0xnorb0 comparator_0/xnor_3/not_0/in vdd comparator_0/xnor_3/not_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1445 comparator_0/a0xnorb0 comparator_0/xnor_3/not_0/in gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1446 comparator_0/xnor_3/not_0/in boout_2 comparator_0/xnor_3/XOR_0/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1447 comparator_0/xnor_3/XOR_0/bbar boout_2 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1448 comparator_0/xnor_3/not_0/in comparator_0/xnor_3/XOR_0/bbar comparator_0/xnor_3/XOR_0/abar comparator_0/xnor_3/XOR_0/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1449 vdd boout_2 comparator_0/xnor_3/XOR_0/bbar comparator_0/xnor_3/XOR_0/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1450 comparator_0/xnor_3/not_0/in boout_2 a0out_2 comparator_0/xnor_3/XOR_0/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1451 comparator_0/xnor_3/XOR_0/abar a0out_2 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1452 vdd a0out_2 comparator_0/xnor_3/XOR_0/abar comparator_0/xnor_3/XOR_0/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1453 comparator_0/xnor_3/not_0/in comparator_0/xnor_3/XOR_0/bbar a0out_2 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1454 comparator_0/a1bar a1out_2 vdd comparator_0/not_5/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1455 comparator_0/a1bar a1out_2 gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1456 comparator_0/a2bar a2out_2 vdd comparator_0/not_6/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1457 comparator_0/a2bar a2out_2 gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1458 comparator_0/a3bar a3out_2 vdd comparator_0/not_7/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1459 comparator_0/a3bar a3out_2 gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1460 comparator_0/t8 comparator_0/5input_AND_0/not_0/in vdd comparator_0/5input_AND_0/not_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1461 comparator_0/t8 comparator_0/5input_AND_0/not_0/in gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1462 vdd a0out_2 comparator_0/5input_AND_0/not_0/in comparator_0/5input_AND_0/w_n37_15# CMOSP w=14 l=8
+  ad=0 pd=0 as=405 ps=198
M1463 vdd comparator_0/a3xnorb3 comparator_0/5input_AND_0/not_0/in comparator_0/5input_AND_0/w_31_n55# CMOSP w=15 l=8
+  ad=0 pd=0 as=0 ps=0
M1464 comparator_0/5input_AND_0/a_n33_n203# comparator_0/b0bar comparator_0/5input_AND_0/a_n33_n226# Gnd CMOSN w=36 l=12
+  ad=468 pd=98 as=396 ps=94
M1465 comparator_0/5input_AND_0/not_0/in comparator_0/a1xnorb1 comparator_0/5input_AND_0/a_n33_n154# Gnd CMOSN w=36 l=12
+  ad=540 pd=102 as=432 ps=96
M1466 vdd comparator_0/a1xnorb1 comparator_0/5input_AND_0/not_0/in comparator_0/5input_AND_0/w_106_n113# CMOSP w=13 l=8
+  ad=0 pd=0 as=0 ps=0
M1467 comparator_0/5input_AND_0/a_n33_n154# comparator_0/a2xnorb2 comparator_0/5input_AND_0/a_n33_n178# Gnd CMOSN w=36 l=12
+  ad=0 pd=0 as=432 ps=96
M1468 comparator_0/5input_AND_0/a_n33_n178# comparator_0/a3xnorb3 comparator_0/5input_AND_0/a_n33_n203# Gnd CMOSN w=36 l=12
+  ad=0 pd=0 as=0 ps=0
M1469 comparator_0/5input_AND_0/a_n33_n226# a0out_2 gnd Gnd CMOSN w=36 l=12
+  ad=0 pd=0 as=0 ps=0
M1470 vdd comparator_0/b0bar comparator_0/5input_AND_0/not_0/in comparator_0/5input_AND_0/w_n4_n20# CMOSP w=13 l=8
+  ad=0 pd=0 as=0 ps=0
M1471 vdd comparator_0/a2xnorb2 comparator_0/5input_AND_0/not_0/in comparator_0/5input_AND_0/w_68_n82# CMOSP w=14 l=8
+  ad=0 pd=0 as=0 ps=0
M1472 comparator_0/t4 comparator_0/5input_AND_1/not_0/in vdd comparator_0/5input_AND_1/not_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1473 comparator_0/t4 comparator_0/5input_AND_1/not_0/in gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1474 vdd comparator_0/a0bar comparator_0/5input_AND_1/not_0/in comparator_0/5input_AND_1/w_n37_15# CMOSP w=14 l=8
+  ad=0 pd=0 as=405 ps=198
M1475 vdd comparator_0/a1xnorb1 comparator_0/5input_AND_1/not_0/in comparator_0/5input_AND_1/w_31_n55# CMOSP w=15 l=8
+  ad=0 pd=0 as=0 ps=0
M1476 comparator_0/5input_AND_1/a_n33_n203# boout_2 comparator_0/5input_AND_1/a_n33_n226# Gnd CMOSN w=36 l=12
+  ad=468 pd=98 as=396 ps=94
M1477 comparator_0/5input_AND_1/not_0/in comparator_0/a3xnorb3 comparator_0/5input_AND_1/a_n33_n154# Gnd CMOSN w=36 l=12
+  ad=540 pd=102 as=432 ps=96
M1478 vdd comparator_0/a3xnorb3 comparator_0/5input_AND_1/not_0/in comparator_0/5input_AND_1/w_106_n113# CMOSP w=13 l=8
+  ad=0 pd=0 as=0 ps=0
M1479 comparator_0/5input_AND_1/a_n33_n154# comparator_0/a2xnorb2 comparator_0/5input_AND_1/a_n33_n178# Gnd CMOSN w=36 l=12
+  ad=0 pd=0 as=432 ps=96
M1480 comparator_0/5input_AND_1/a_n33_n178# comparator_0/a1xnorb1 comparator_0/5input_AND_1/a_n33_n203# Gnd CMOSN w=36 l=12
+  ad=0 pd=0 as=0 ps=0
M1481 comparator_0/5input_AND_1/a_n33_n226# comparator_0/a0bar gnd Gnd CMOSN w=36 l=12
+  ad=0 pd=0 as=0 ps=0
M1482 vdd boout_2 comparator_0/5input_AND_1/not_0/in comparator_0/5input_AND_1/w_n4_n20# CMOSP w=13 l=8
+  ad=0 pd=0 as=0 ps=0
M1483 vdd comparator_0/a2xnorb2 comparator_0/5input_AND_1/not_0/in comparator_0/5input_AND_1/w_68_n82# CMOSP w=14 l=8
+  ad=0 pd=0 as=0 ps=0
M1484 comparator_0/t5 comparator_0/and_0/a_n26_14# vdd comparator_0/and_0/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1485 vdd comparator_0/b3bar comparator_0/and_0/a_n26_14# comparator_0/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1486 comparator_0/t5 comparator_0/and_0/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1487 comparator_0/and_0/a_n26_14# a3out_2 vdd comparator_0/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1488 comparator_0/and_0/a_n26_n23# a3out_2 gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1489 comparator_0/and_0/a_n26_14# comparator_0/b3bar comparator_0/and_0/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1490 equal comparator_0/4input_AND_0/not_0/in vdd comparator_0/4input_AND_0/not_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1491 equal comparator_0/4input_AND_0/not_0/in gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1492 vdd comparator_0/a3xnorb3 comparator_0/4input_AND_0/not_0/in comparator_0/4input_AND_0/w_n47_52# CMOSP w=12 l=7
+  ad=0 pd=0 as=648 ps=204
M1493 comparator_0/4input_AND_0/not_0/in comparator_0/a0xnorb0 comparator_0/4input_AND_0/a_n40_n132# Gnd CMOSN w=12 l=7
+  ad=120 pd=44 as=96 ps=40
M1494 comparator_0/4input_AND_0/a_n40_n147# comparator_0/a2xnorb2 comparator_0/4input_AND_0/a_n40_n162# Gnd CMOSN w=12 l=7
+  ad=96 pd=40 as=96 ps=40
M1495 vdd comparator_0/a0xnorb0 comparator_0/4input_AND_0/not_0/in comparator_0/4input_AND_0/w_68_n95# CMOSP w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1496 comparator_0/4input_AND_0/a_n40_n132# comparator_0/a1xnorb1 comparator_0/4input_AND_0/a_n40_n147# Gnd CMOSN w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1497 comparator_0/4input_AND_0/a_n40_n162# comparator_0/a3xnorb3 gnd Gnd CMOSN w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1498 vdd comparator_0/a2xnorb2 comparator_0/4input_AND_0/not_0/in comparator_0/4input_AND_0/w_n8_2# CMOSP w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1499 vdd comparator_0/a1xnorb1 comparator_0/4input_AND_0/not_0/in comparator_0/4input_AND_0/w_29_n46# CMOSP w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1500 comparator_0/t7 comparator_0/4input_AND_1/not_0/in vdd comparator_0/4input_AND_1/not_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1501 comparator_0/t7 comparator_0/4input_AND_1/not_0/in gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1502 vdd a1out_2 comparator_0/4input_AND_1/not_0/in comparator_0/4input_AND_1/w_n47_52# CMOSP w=12 l=7
+  ad=0 pd=0 as=648 ps=204
M1503 comparator_0/4input_AND_1/not_0/in comparator_0/a2xnorb2 comparator_0/4input_AND_1/a_n40_n132# Gnd CMOSN w=12 l=7
+  ad=120 pd=44 as=96 ps=40
M1504 comparator_0/4input_AND_1/a_n40_n147# comparator_0/b1bar comparator_0/4input_AND_1/a_n40_n162# Gnd CMOSN w=12 l=7
+  ad=96 pd=40 as=96 ps=40
M1505 vdd comparator_0/a2xnorb2 comparator_0/4input_AND_1/not_0/in comparator_0/4input_AND_1/w_68_n95# CMOSP w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1506 comparator_0/4input_AND_1/a_n40_n132# comparator_0/a3xnorb3 comparator_0/4input_AND_1/a_n40_n147# Gnd CMOSN w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1507 comparator_0/4input_AND_1/a_n40_n162# a1out_2 gnd Gnd CMOSN w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1508 vdd comparator_0/b1bar comparator_0/4input_AND_1/not_0/in comparator_0/4input_AND_1/w_n8_2# CMOSP w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1509 vdd comparator_0/a3xnorb3 comparator_0/4input_AND_1/not_0/in comparator_0/4input_AND_1/w_29_n46# CMOSP w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1510 comparator_0/t1 comparator_0/and_1/a_n26_14# vdd comparator_0/and_1/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1511 vdd comparator_0/b3 comparator_0/and_1/a_n26_14# comparator_0/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1512 comparator_0/t1 comparator_0/and_1/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1513 comparator_0/and_1/a_n26_14# comparator_0/a3bar vdd comparator_0/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1514 comparator_0/and_1/a_n26_n23# comparator_0/a3bar gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1515 comparator_0/and_1/a_n26_14# comparator_0/b3 comparator_0/and_1/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1516 comparator_0/t3 comparator_0/4input_AND_2/not_0/in vdd comparator_0/4input_AND_2/not_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1517 comparator_0/t3 comparator_0/4input_AND_2/not_0/in gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1518 vdd comparator_0/a1bar comparator_0/4input_AND_2/not_0/in comparator_0/4input_AND_2/w_n47_52# CMOSP w=12 l=7
+  ad=0 pd=0 as=648 ps=204
M1519 comparator_0/4input_AND_2/not_0/in comparator_0/a3xnorb3 comparator_0/4input_AND_2/a_n40_n132# Gnd CMOSN w=12 l=7
+  ad=120 pd=44 as=96 ps=40
M1520 comparator_0/4input_AND_2/a_n40_n147# b1out_2 comparator_0/4input_AND_2/a_n40_n162# Gnd CMOSN w=12 l=7
+  ad=96 pd=40 as=96 ps=40
M1521 vdd comparator_0/a3xnorb3 comparator_0/4input_AND_2/not_0/in comparator_0/4input_AND_2/w_68_n95# CMOSP w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1522 comparator_0/4input_AND_2/a_n40_n132# comparator_0/a2xnorb2 comparator_0/4input_AND_2/a_n40_n147# Gnd CMOSN w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1523 comparator_0/4input_AND_2/a_n40_n162# comparator_0/a1bar gnd Gnd CMOSN w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1524 vdd b1out_2 comparator_0/4input_AND_2/not_0/in comparator_0/4input_AND_2/w_n8_2# CMOSP w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1525 vdd comparator_0/a2xnorb2 comparator_0/4input_AND_2/not_0/in comparator_0/4input_AND_2/w_29_n46# CMOSP w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1526 comparator_0/t6 comparator_0/3input_AND_0/not_0/in vdd comparator_0/3input_AND_0/not_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1527 comparator_0/t6 comparator_0/3input_AND_0/not_0/in gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1528 comparator_0/3input_AND_0/a_n9_n125# comparator_0/b2bar gnd Gnd CMOSN w=15 l=8
+  ad=135 pd=48 as=0 ps=0
M1529 comparator_0/3input_AND_0/not_0/in comparator_0/a3xnorb3 comparator_0/3input_AND_0/a_n9_n108# Gnd CMOSN w=15 l=8
+  ad=165 pd=52 as=165 ps=52
M1530 vdd comparator_0/a3xnorb3 comparator_0/3input_AND_0/not_0/in comparator_0/3input_AND_0/w_69_n71# CMOSP w=13 l=8
+  ad=0 pd=0 as=546 ps=162
M1531 vdd a2out_2 comparator_0/3input_AND_0/not_0/in comparator_0/3input_AND_0/w_32_n21# CMOSP w=13 l=8
+  ad=0 pd=0 as=0 ps=0
M1532 vdd comparator_0/b2bar comparator_0/3input_AND_0/not_0/in comparator_0/3input_AND_0/w_n14_24# CMOSP w=13 l=8
+  ad=0 pd=0 as=0 ps=0
M1533 comparator_0/3input_AND_0/a_n9_n108# a2out_2 comparator_0/3input_AND_0/a_n9_n125# Gnd CMOSN w=15 l=8
+  ad=0 pd=0 as=0 ps=0
M1534 comparator_0/t2 comparator_0/3input_AND_1/not_0/in vdd comparator_0/3input_AND_1/not_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1535 comparator_0/t2 comparator_0/3input_AND_1/not_0/in gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1536 comparator_0/3input_AND_1/a_n9_n125# comparator_0/a2bar gnd Gnd CMOSN w=15 l=8
+  ad=135 pd=48 as=0 ps=0
M1537 comparator_0/3input_AND_1/not_0/in comparator_0/a3xnorb3 comparator_0/3input_AND_1/a_n9_n108# Gnd CMOSN w=15 l=8
+  ad=165 pd=52 as=165 ps=52
M1538 vdd comparator_0/a3xnorb3 comparator_0/3input_AND_1/not_0/in comparator_0/3input_AND_1/w_69_n71# CMOSP w=13 l=8
+  ad=0 pd=0 as=546 ps=162
M1539 vdd b2out_2 comparator_0/3input_AND_1/not_0/in comparator_0/3input_AND_1/w_32_n21# CMOSP w=13 l=8
+  ad=0 pd=0 as=0 ps=0
M1540 vdd comparator_0/a2bar comparator_0/3input_AND_1/not_0/in comparator_0/3input_AND_1/w_n14_24# CMOSP w=13 l=8
+  ad=0 pd=0 as=0 ps=0
M1541 comparator_0/3input_AND_1/a_n9_n108# b2out_2 comparator_0/3input_AND_1/a_n9_n125# Gnd CMOSN w=15 l=8
+  ad=0 pd=0 as=0 ps=0
M1542 4bitadder_1/fulladder_0/or_0/a_n15_32# 4bitadder_1/fulladder_0/or_0/a gnd Gnd CMOSN w=16 l=5
+  ad=304 pd=70 as=0 ps=0
M1543 4bitadder_1/c1 4bitadder_1/fulladder_0/or_0/a_n15_32# vdd 4bitadder_1/fulladder_0/or_0/w_58_101# CMOSP w=16 l=6
+  ad=288 pd=68 as=0 ps=0
M1544 gnd 4bitadder_1/fulladder_0/or_0/b 4bitadder_1/fulladder_0/or_0/a_n15_32# Gnd CMOSN w=16 l=5
+  ad=0 pd=0 as=0 ps=0
M1545 4bitadder_1/fulladder_0/or_0/a_n15_32# 4bitadder_1/fulladder_0/or_0/b 4bitadder_1/fulladder_0/or_0/a_n15_107# 4bitadder_1/fulladder_0/or_0/w_n48_101# CMOSP w=16 l=5
+  ad=448 pd=88 as=304 ps=70
M1546 4bitadder_1/c1 4bitadder_1/fulladder_0/or_0/a_n15_32# gnd Gnd CMOSN w=16 l=6
+  ad=320 pd=72 as=0 ps=0
M1547 4bitadder_1/fulladder_0/or_0/a_n15_107# 4bitadder_1/fulladder_0/or_0/a vdd 4bitadder_1/fulladder_0/or_0/w_n48_101# CMOSP w=16 l=5
+  ad=0 pd=0 as=0 ps=0
M1548 4bitadder_1/fulladder_0/or_0/a 4bitadder_1/fulladder_0/and_0/a_n26_14# vdd 4bitadder_1/fulladder_0/and_0/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1549 vdd s0 4bitadder_1/fulladder_0/and_0/a_n26_14# 4bitadder_1/fulladder_0/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1550 4bitadder_1/fulladder_0/or_0/a 4bitadder_1/fulladder_0/and_0/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1551 4bitadder_1/fulladder_0/and_0/a_n26_14# 4bitadder_1/fulladder_0/axorb vdd 4bitadder_1/fulladder_0/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1552 4bitadder_1/fulladder_0/and_0/a_n26_n23# 4bitadder_1/fulladder_0/axorb gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1553 4bitadder_1/fulladder_0/and_0/a_n26_14# s0 4bitadder_1/fulladder_0/and_0/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1554 4bitadder_1/fulladder_0/axorb 4bitadder_1/b0xorM 4bitadder_1/fulladder_0/XOR_0/abar Gnd CMOSN w=11 l=6
+  ad=495 pd=156 as=407 ps=118
M1555 4bitadder_1/fulladder_0/XOR_0/bbar 4bitadder_1/b0xorM gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1556 4bitadder_1/fulladder_0/axorb 4bitadder_1/fulladder_0/XOR_0/bbar 4bitadder_1/fulladder_0/XOR_0/abar 4bitadder_1/fulladder_0/XOR_0/w_62_n20# CMOSP w=12 l=6
+  ad=252 pd=110 as=218 ps=84
M1557 vdd 4bitadder_1/b0xorM 4bitadder_1/fulladder_0/XOR_0/bbar 4bitadder_1/fulladder_0/XOR_0/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1558 4bitadder_1/fulladder_0/axorb 4bitadder_1/b0xorM a0_out1 4bitadder_1/fulladder_0/XOR_0/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1559 4bitadder_1/fulladder_0/XOR_0/abar a0_out1 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1560 vdd a0_out1 4bitadder_1/fulladder_0/XOR_0/abar 4bitadder_1/fulladder_0/XOR_0/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1561 4bitadder_1/fulladder_0/axorb 4bitadder_1/fulladder_0/XOR_0/bbar a0_out1 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1562 4bitadder_1/fulladder_0/or_0/b 4bitadder_1/fulladder_0/and_1/a_n26_14# vdd 4bitadder_1/fulladder_0/and_1/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1563 vdd a0_out1 4bitadder_1/fulladder_0/and_1/a_n26_14# 4bitadder_1/fulladder_0/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1564 4bitadder_1/fulladder_0/or_0/b 4bitadder_1/fulladder_0/and_1/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1565 4bitadder_1/fulladder_0/and_1/a_n26_14# 4bitadder_1/b0xorM vdd 4bitadder_1/fulladder_0/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1566 4bitadder_1/fulladder_0/and_1/a_n26_n23# 4bitadder_1/b0xorM gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1567 4bitadder_1/fulladder_0/and_1/a_n26_14# a0_out1 4bitadder_1/fulladder_0/and_1/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1568 s0_sub s0 4bitadder_1/fulladder_0/XOR_1/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1569 4bitadder_1/fulladder_0/XOR_1/bbar s0 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1570 s0_sub 4bitadder_1/fulladder_0/XOR_1/bbar 4bitadder_1/fulladder_0/XOR_1/abar 4bitadder_1/fulladder_0/XOR_1/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1571 vdd s0 4bitadder_1/fulladder_0/XOR_1/bbar 4bitadder_1/fulladder_0/XOR_1/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1572 s0_sub s0 4bitadder_1/fulladder_0/axorb 4bitadder_1/fulladder_0/XOR_1/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1573 4bitadder_1/fulladder_0/XOR_1/abar 4bitadder_1/fulladder_0/axorb gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1574 vdd 4bitadder_1/fulladder_0/axorb 4bitadder_1/fulladder_0/XOR_1/abar 4bitadder_1/fulladder_0/XOR_1/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1575 s0_sub 4bitadder_1/fulladder_0/XOR_1/bbar 4bitadder_1/fulladder_0/axorb Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1576 4bitadder_1/fulladder_1/or_0/a_n15_32# 4bitadder_1/fulladder_1/or_0/a gnd Gnd CMOSN w=16 l=5
+  ad=304 pd=70 as=0 ps=0
M1577 4bitadder_1/c2 4bitadder_1/fulladder_1/or_0/a_n15_32# vdd 4bitadder_1/fulladder_1/or_0/w_58_101# CMOSP w=16 l=6
+  ad=288 pd=68 as=0 ps=0
M1578 gnd 4bitadder_1/fulladder_1/or_0/b 4bitadder_1/fulladder_1/or_0/a_n15_32# Gnd CMOSN w=16 l=5
+  ad=0 pd=0 as=0 ps=0
M1579 4bitadder_1/fulladder_1/or_0/a_n15_32# 4bitadder_1/fulladder_1/or_0/b 4bitadder_1/fulladder_1/or_0/a_n15_107# 4bitadder_1/fulladder_1/or_0/w_n48_101# CMOSP w=16 l=5
+  ad=448 pd=88 as=304 ps=70
M1580 4bitadder_1/c2 4bitadder_1/fulladder_1/or_0/a_n15_32# gnd Gnd CMOSN w=16 l=6
+  ad=320 pd=72 as=0 ps=0
M1581 4bitadder_1/fulladder_1/or_0/a_n15_107# 4bitadder_1/fulladder_1/or_0/a vdd 4bitadder_1/fulladder_1/or_0/w_n48_101# CMOSP w=16 l=5
+  ad=0 pd=0 as=0 ps=0
M1582 4bitadder_1/fulladder_1/or_0/a 4bitadder_1/fulladder_1/and_0/a_n26_14# vdd 4bitadder_1/fulladder_1/and_0/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1583 vdd 4bitadder_1/c1 4bitadder_1/fulladder_1/and_0/a_n26_14# 4bitadder_1/fulladder_1/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1584 4bitadder_1/fulladder_1/or_0/a 4bitadder_1/fulladder_1/and_0/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1585 4bitadder_1/fulladder_1/and_0/a_n26_14# 4bitadder_1/fulladder_1/axorb vdd 4bitadder_1/fulladder_1/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1586 4bitadder_1/fulladder_1/and_0/a_n26_n23# 4bitadder_1/fulladder_1/axorb gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1587 4bitadder_1/fulladder_1/and_0/a_n26_14# 4bitadder_1/c1 4bitadder_1/fulladder_1/and_0/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1588 4bitadder_1/fulladder_1/axorb 4bitadder_1/XOR_1/out 4bitadder_1/fulladder_1/XOR_0/abar Gnd CMOSN w=11 l=6
+  ad=495 pd=156 as=407 ps=118
M1589 4bitadder_1/fulladder_1/XOR_0/bbar 4bitadder_1/XOR_1/out gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1590 4bitadder_1/fulladder_1/axorb 4bitadder_1/fulladder_1/XOR_0/bbar 4bitadder_1/fulladder_1/XOR_0/abar 4bitadder_1/fulladder_1/XOR_0/w_62_n20# CMOSP w=12 l=6
+  ad=252 pd=110 as=218 ps=84
M1591 vdd 4bitadder_1/XOR_1/out 4bitadder_1/fulladder_1/XOR_0/bbar 4bitadder_1/fulladder_1/XOR_0/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1592 4bitadder_1/fulladder_1/axorb 4bitadder_1/XOR_1/out a1out_1 4bitadder_1/fulladder_1/XOR_0/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1593 4bitadder_1/fulladder_1/XOR_0/abar a1out_1 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1594 vdd a1out_1 4bitadder_1/fulladder_1/XOR_0/abar 4bitadder_1/fulladder_1/XOR_0/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1595 4bitadder_1/fulladder_1/axorb 4bitadder_1/fulladder_1/XOR_0/bbar a1out_1 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1596 4bitadder_1/fulladder_1/or_0/b 4bitadder_1/fulladder_1/and_1/a_n26_14# vdd 4bitadder_1/fulladder_1/and_1/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1597 vdd a1out_1 4bitadder_1/fulladder_1/and_1/a_n26_14# 4bitadder_1/fulladder_1/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1598 4bitadder_1/fulladder_1/or_0/b 4bitadder_1/fulladder_1/and_1/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1599 4bitadder_1/fulladder_1/and_1/a_n26_14# 4bitadder_1/XOR_1/out vdd 4bitadder_1/fulladder_1/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1600 4bitadder_1/fulladder_1/and_1/a_n26_n23# 4bitadder_1/XOR_1/out gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1601 4bitadder_1/fulladder_1/and_1/a_n26_14# a1out_1 4bitadder_1/fulladder_1/and_1/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1602 s1_sub 4bitadder_1/c1 4bitadder_1/fulladder_1/XOR_1/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1603 4bitadder_1/fulladder_1/XOR_1/bbar 4bitadder_1/c1 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1604 s1_sub 4bitadder_1/fulladder_1/XOR_1/bbar 4bitadder_1/fulladder_1/XOR_1/abar 4bitadder_1/fulladder_1/XOR_1/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1605 vdd 4bitadder_1/c1 4bitadder_1/fulladder_1/XOR_1/bbar 4bitadder_1/fulladder_1/XOR_1/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1606 s1_sub 4bitadder_1/c1 4bitadder_1/fulladder_1/axorb 4bitadder_1/fulladder_1/XOR_1/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1607 4bitadder_1/fulladder_1/XOR_1/abar 4bitadder_1/fulladder_1/axorb gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1608 vdd 4bitadder_1/fulladder_1/axorb 4bitadder_1/fulladder_1/XOR_1/abar 4bitadder_1/fulladder_1/XOR_1/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1609 s1_sub 4bitadder_1/fulladder_1/XOR_1/bbar 4bitadder_1/fulladder_1/axorb Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1610 4bitadder_1/fulladder_2/or_0/a_n15_32# 4bitadder_1/fulladder_2/or_0/a gnd Gnd CMOSN w=16 l=5
+  ad=304 pd=70 as=0 ps=0
M1611 4bitadder_1/c3 4bitadder_1/fulladder_2/or_0/a_n15_32# vdd 4bitadder_1/fulladder_2/or_0/w_58_101# CMOSP w=16 l=6
+  ad=288 pd=68 as=0 ps=0
M1612 gnd 4bitadder_1/fulladder_2/or_0/b 4bitadder_1/fulladder_2/or_0/a_n15_32# Gnd CMOSN w=16 l=5
+  ad=0 pd=0 as=0 ps=0
M1613 4bitadder_1/fulladder_2/or_0/a_n15_32# 4bitadder_1/fulladder_2/or_0/b 4bitadder_1/fulladder_2/or_0/a_n15_107# 4bitadder_1/fulladder_2/or_0/w_n48_101# CMOSP w=16 l=5
+  ad=448 pd=88 as=304 ps=70
M1614 4bitadder_1/c3 4bitadder_1/fulladder_2/or_0/a_n15_32# gnd Gnd CMOSN w=16 l=6
+  ad=320 pd=72 as=0 ps=0
M1615 4bitadder_1/fulladder_2/or_0/a_n15_107# 4bitadder_1/fulladder_2/or_0/a vdd 4bitadder_1/fulladder_2/or_0/w_n48_101# CMOSP w=16 l=5
+  ad=0 pd=0 as=0 ps=0
M1616 4bitadder_1/fulladder_2/or_0/a 4bitadder_1/fulladder_2/and_0/a_n26_14# vdd 4bitadder_1/fulladder_2/and_0/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1617 vdd 4bitadder_1/c2 4bitadder_1/fulladder_2/and_0/a_n26_14# 4bitadder_1/fulladder_2/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1618 4bitadder_1/fulladder_2/or_0/a 4bitadder_1/fulladder_2/and_0/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1619 4bitadder_1/fulladder_2/and_0/a_n26_14# 4bitadder_1/fulladder_2/axorb vdd 4bitadder_1/fulladder_2/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1620 4bitadder_1/fulladder_2/and_0/a_n26_n23# 4bitadder_1/fulladder_2/axorb gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1621 4bitadder_1/fulladder_2/and_0/a_n26_14# 4bitadder_1/c2 4bitadder_1/fulladder_2/and_0/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1622 4bitadder_1/fulladder_2/axorb 4bitadder_1/XOR_2/out 4bitadder_1/fulladder_2/XOR_0/abar Gnd CMOSN w=11 l=6
+  ad=495 pd=156 as=407 ps=118
M1623 4bitadder_1/fulladder_2/XOR_0/bbar 4bitadder_1/XOR_2/out gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1624 4bitadder_1/fulladder_2/axorb 4bitadder_1/fulladder_2/XOR_0/bbar 4bitadder_1/fulladder_2/XOR_0/abar 4bitadder_1/fulladder_2/XOR_0/w_62_n20# CMOSP w=12 l=6
+  ad=252 pd=110 as=218 ps=84
M1625 vdd 4bitadder_1/XOR_2/out 4bitadder_1/fulladder_2/XOR_0/bbar 4bitadder_1/fulladder_2/XOR_0/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1626 4bitadder_1/fulladder_2/axorb 4bitadder_1/XOR_2/out a2out_1 4bitadder_1/fulladder_2/XOR_0/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1627 4bitadder_1/fulladder_2/XOR_0/abar a2out_1 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1628 vdd a2out_1 4bitadder_1/fulladder_2/XOR_0/abar 4bitadder_1/fulladder_2/XOR_0/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1629 4bitadder_1/fulladder_2/axorb 4bitadder_1/fulladder_2/XOR_0/bbar a2out_1 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1630 4bitadder_1/fulladder_2/or_0/b 4bitadder_1/fulladder_2/and_1/a_n26_14# vdd 4bitadder_1/fulladder_2/and_1/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1631 vdd a2out_1 4bitadder_1/fulladder_2/and_1/a_n26_14# 4bitadder_1/fulladder_2/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1632 4bitadder_1/fulladder_2/or_0/b 4bitadder_1/fulladder_2/and_1/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1633 4bitadder_1/fulladder_2/and_1/a_n26_14# 4bitadder_1/XOR_2/out vdd 4bitadder_1/fulladder_2/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1634 4bitadder_1/fulladder_2/and_1/a_n26_n23# 4bitadder_1/XOR_2/out gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1635 4bitadder_1/fulladder_2/and_1/a_n26_14# a2out_1 4bitadder_1/fulladder_2/and_1/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1636 s2_sub 4bitadder_1/c2 4bitadder_1/fulladder_2/XOR_1/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1637 4bitadder_1/fulladder_2/XOR_1/bbar 4bitadder_1/c2 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1638 s2_sub 4bitadder_1/fulladder_2/XOR_1/bbar 4bitadder_1/fulladder_2/XOR_1/abar 4bitadder_1/fulladder_2/XOR_1/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1639 vdd 4bitadder_1/c2 4bitadder_1/fulladder_2/XOR_1/bbar 4bitadder_1/fulladder_2/XOR_1/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1640 s2_sub 4bitadder_1/c2 4bitadder_1/fulladder_2/axorb 4bitadder_1/fulladder_2/XOR_1/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1641 4bitadder_1/fulladder_2/XOR_1/abar 4bitadder_1/fulladder_2/axorb gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1642 vdd 4bitadder_1/fulladder_2/axorb 4bitadder_1/fulladder_2/XOR_1/abar 4bitadder_1/fulladder_2/XOR_1/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1643 s2_sub 4bitadder_1/fulladder_2/XOR_1/bbar 4bitadder_1/fulladder_2/axorb Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1644 4bitadder_1/fulladder_3/or_0/a_n15_32# 4bitadder_1/fulladder_3/or_0/a gnd Gnd CMOSN w=16 l=5
+  ad=304 pd=70 as=0 ps=0
M1645 fc_sub 4bitadder_1/fulladder_3/or_0/a_n15_32# vdd 4bitadder_1/fulladder_3/or_0/w_58_101# CMOSP w=16 l=6
+  ad=288 pd=68 as=0 ps=0
M1646 gnd 4bitadder_1/fulladder_3/or_0/b 4bitadder_1/fulladder_3/or_0/a_n15_32# Gnd CMOSN w=16 l=5
+  ad=0 pd=0 as=0 ps=0
M1647 4bitadder_1/fulladder_3/or_0/a_n15_32# 4bitadder_1/fulladder_3/or_0/b 4bitadder_1/fulladder_3/or_0/a_n15_107# 4bitadder_1/fulladder_3/or_0/w_n48_101# CMOSP w=16 l=5
+  ad=448 pd=88 as=304 ps=70
M1648 fc_sub 4bitadder_1/fulladder_3/or_0/a_n15_32# gnd Gnd CMOSN w=16 l=6
+  ad=320 pd=72 as=0 ps=0
M1649 4bitadder_1/fulladder_3/or_0/a_n15_107# 4bitadder_1/fulladder_3/or_0/a vdd 4bitadder_1/fulladder_3/or_0/w_n48_101# CMOSP w=16 l=5
+  ad=0 pd=0 as=0 ps=0
M1650 4bitadder_1/fulladder_3/or_0/a 4bitadder_1/fulladder_3/and_0/a_n26_14# vdd 4bitadder_1/fulladder_3/and_0/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1651 vdd 4bitadder_1/c3 4bitadder_1/fulladder_3/and_0/a_n26_14# 4bitadder_1/fulladder_3/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1652 4bitadder_1/fulladder_3/or_0/a 4bitadder_1/fulladder_3/and_0/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1653 4bitadder_1/fulladder_3/and_0/a_n26_14# 4bitadder_1/fulladder_3/axorb vdd 4bitadder_1/fulladder_3/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1654 4bitadder_1/fulladder_3/and_0/a_n26_n23# 4bitadder_1/fulladder_3/axorb gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1655 4bitadder_1/fulladder_3/and_0/a_n26_14# 4bitadder_1/c3 4bitadder_1/fulladder_3/and_0/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1656 4bitadder_1/fulladder_3/axorb 4bitadder_1/XOR_3/out 4bitadder_1/fulladder_3/XOR_0/abar Gnd CMOSN w=11 l=6
+  ad=495 pd=156 as=407 ps=118
M1657 4bitadder_1/fulladder_3/XOR_0/bbar 4bitadder_1/XOR_3/out gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1658 4bitadder_1/fulladder_3/axorb 4bitadder_1/fulladder_3/XOR_0/bbar 4bitadder_1/fulladder_3/XOR_0/abar 4bitadder_1/fulladder_3/XOR_0/w_62_n20# CMOSP w=12 l=6
+  ad=252 pd=110 as=218 ps=84
M1659 vdd 4bitadder_1/XOR_3/out 4bitadder_1/fulladder_3/XOR_0/bbar 4bitadder_1/fulladder_3/XOR_0/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1660 4bitadder_1/fulladder_3/axorb 4bitadder_1/XOR_3/out a3out_1 4bitadder_1/fulladder_3/XOR_0/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1661 4bitadder_1/fulladder_3/XOR_0/abar a3out_1 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1662 vdd a3out_1 4bitadder_1/fulladder_3/XOR_0/abar 4bitadder_1/fulladder_3/XOR_0/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1663 4bitadder_1/fulladder_3/axorb 4bitadder_1/fulladder_3/XOR_0/bbar a3out_1 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1664 4bitadder_1/fulladder_3/or_0/b 4bitadder_1/fulladder_3/and_1/a_n26_14# vdd 4bitadder_1/fulladder_3/and_1/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1665 vdd a3out_1 4bitadder_1/fulladder_3/and_1/a_n26_14# 4bitadder_1/fulladder_3/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1666 4bitadder_1/fulladder_3/or_0/b 4bitadder_1/fulladder_3/and_1/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1667 4bitadder_1/fulladder_3/and_1/a_n26_14# 4bitadder_1/XOR_3/out vdd 4bitadder_1/fulladder_3/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1668 4bitadder_1/fulladder_3/and_1/a_n26_n23# 4bitadder_1/XOR_3/out gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1669 4bitadder_1/fulladder_3/and_1/a_n26_14# a3out_1 4bitadder_1/fulladder_3/and_1/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1670 s3_sub 4bitadder_1/c3 4bitadder_1/fulladder_3/XOR_1/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1671 4bitadder_1/fulladder_3/XOR_1/bbar 4bitadder_1/c3 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1672 s3_sub 4bitadder_1/fulladder_3/XOR_1/bbar 4bitadder_1/fulladder_3/XOR_1/abar 4bitadder_1/fulladder_3/XOR_1/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1673 vdd 4bitadder_1/c3 4bitadder_1/fulladder_3/XOR_1/bbar 4bitadder_1/fulladder_3/XOR_1/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1674 s3_sub 4bitadder_1/c3 4bitadder_1/fulladder_3/axorb 4bitadder_1/fulladder_3/XOR_1/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1675 4bitadder_1/fulladder_3/XOR_1/abar 4bitadder_1/fulladder_3/axorb gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1676 vdd 4bitadder_1/fulladder_3/axorb 4bitadder_1/fulladder_3/XOR_1/abar 4bitadder_1/fulladder_3/XOR_1/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1677 s3_sub 4bitadder_1/fulladder_3/XOR_1/bbar 4bitadder_1/fulladder_3/axorb Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1678 4bitadder_1/b0xorM s0 4bitadder_1/XOR_0/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1679 4bitadder_1/XOR_0/bbar s0 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1680 4bitadder_1/b0xorM 4bitadder_1/XOR_0/bbar 4bitadder_1/XOR_0/abar 4bitadder_1/XOR_0/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1681 vdd s0 4bitadder_1/XOR_0/bbar 4bitadder_1/XOR_0/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1682 4bitadder_1/b0xorM s0 b0out_1 4bitadder_1/XOR_0/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1683 4bitadder_1/XOR_0/abar b0out_1 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1684 vdd b0out_1 4bitadder_1/XOR_0/abar 4bitadder_1/XOR_0/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1685 4bitadder_1/b0xorM 4bitadder_1/XOR_0/bbar b0out_1 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1686 4bitadder_1/XOR_1/out s0 4bitadder_1/XOR_1/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1687 4bitadder_1/XOR_1/bbar s0 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1688 4bitadder_1/XOR_1/out 4bitadder_1/XOR_1/bbar 4bitadder_1/XOR_1/abar 4bitadder_1/XOR_1/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1689 vdd s0 4bitadder_1/XOR_1/bbar 4bitadder_1/XOR_1/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1690 4bitadder_1/XOR_1/out s0 b1out_1 4bitadder_1/XOR_1/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1691 4bitadder_1/XOR_1/abar b1out_1 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1692 vdd b1out_1 4bitadder_1/XOR_1/abar 4bitadder_1/XOR_1/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1693 4bitadder_1/XOR_1/out 4bitadder_1/XOR_1/bbar b1out_1 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1694 4bitadder_1/XOR_2/out s0 4bitadder_1/XOR_2/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1695 4bitadder_1/XOR_2/bbar s0 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1696 4bitadder_1/XOR_2/out 4bitadder_1/XOR_2/bbar 4bitadder_1/XOR_2/abar 4bitadder_1/XOR_2/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1697 vdd s0 4bitadder_1/XOR_2/bbar 4bitadder_1/XOR_2/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1698 4bitadder_1/XOR_2/out s0 b2out_1 4bitadder_1/XOR_2/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1699 4bitadder_1/XOR_2/abar b2out_1 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1700 vdd b2out_1 4bitadder_1/XOR_2/abar 4bitadder_1/XOR_2/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1701 4bitadder_1/XOR_2/out 4bitadder_1/XOR_2/bbar b2out_1 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1702 4bitadder_1/XOR_3/out s0 4bitadder_1/XOR_3/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1703 4bitadder_1/XOR_3/bbar s0 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1704 4bitadder_1/XOR_3/out 4bitadder_1/XOR_3/bbar 4bitadder_1/XOR_3/abar 4bitadder_1/XOR_3/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1705 vdd s0 4bitadder_1/XOR_3/bbar 4bitadder_1/XOR_3/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1706 4bitadder_1/XOR_3/out s0 b3out_1 4bitadder_1/XOR_3/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1707 4bitadder_1/XOR_3/abar b3out_1 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1708 vdd b3out_1 4bitadder_1/XOR_3/abar 4bitadder_1/XOR_3/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1709 4bitadder_1/XOR_3/out 4bitadder_1/XOR_3/bbar b3out_1 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1710 decoder_0/and_2/a s0 vdd decoder_0/not_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1711 decoder_0/and_2/a s0 gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1712 decoder_0/and_1/b s1 vdd decoder_0/not_1/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1713 decoder_0/and_1/b s1 gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1714 enable_0/en decoder_0/and_0/a_n26_14# vdd decoder_0/and_0/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1715 vdd decoder_0/and_1/b decoder_0/and_0/a_n26_14# decoder_0/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1716 enable_0/en decoder_0/and_0/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1717 decoder_0/and_0/a_n26_14# decoder_0/and_2/a vdd decoder_0/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1718 decoder_0/and_0/a_n26_n23# decoder_0/and_2/a gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1719 decoder_0/and_0/a_n26_14# decoder_0/and_1/b decoder_0/and_0/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1720 enable_1/en decoder_0/and_1/a_n26_14# vdd decoder_0/and_1/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1721 vdd decoder_0/and_1/b decoder_0/and_1/a_n26_14# decoder_0/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1722 enable_1/en decoder_0/and_1/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1723 decoder_0/and_1/a_n26_14# s0 vdd decoder_0/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1724 decoder_0/and_1/a_n26_n23# s0 gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1725 decoder_0/and_1/a_n26_14# decoder_0/and_1/b decoder_0/and_1/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1726 enable_2/en decoder_0/and_2/a_n26_14# vdd decoder_0/and_2/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1727 vdd s1 decoder_0/and_2/a_n26_14# decoder_0/and_2/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1728 enable_2/en decoder_0/and_2/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1729 decoder_0/and_2/a_n26_14# decoder_0/and_2/a vdd decoder_0/and_2/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1730 decoder_0/and_2/a_n26_n23# decoder_0/and_2/a gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1731 decoder_0/and_2/a_n26_14# s1 decoder_0/and_2/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1732 enable_3/en decoder_0/and_3/a_n26_14# vdd decoder_0/and_3/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1733 vdd s1 decoder_0/and_3/a_n26_14# decoder_0/and_3/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1734 enable_3/en decoder_0/and_3/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1735 decoder_0/and_3/a_n26_14# s0 vdd decoder_0/and_3/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1736 decoder_0/and_3/a_n26_n23# s0 gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1737 decoder_0/and_3/a_n26_14# s1 decoder_0/and_3/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
C0 a1out_1 4bitadder_1/c1 0.36fF
C1 comparator_0/b3bar comparator_0/a3xnorb3 0.14fF
C2 4bitadder_0/fulladder_1/and_0/a_n26_14# 4bitadder_0/c1 0.10fF
C3 comparator_0/4input_AND_2/w_68_n95# comparator_0/a3xnorb3 0.16fF
C4 4bitadder_0/fulladder_2/and_0/w_n43_8# 4bitadder_0/fulladder_2/axorb 0.09fF
C5 enable_0/and_2/w_n43_8# enable_0/and_2/a_n26_14# 0.02fF
C6 4bitadder_1/fulladder_0/XOR_0/bbar 4bitadder_1/fulladder_0/XOR_0/w_16_n1# 0.03fF
C7 comparator_0/a1xnorb1 comparator_0/xnor_2/not_0/w_n2_10# 0.03fF
C8 4bitadder_1/fulladder_3/XOR_0/w_n34_n1# 4bitadder_1/fulladder_3/XOR_0/abar 0.03fF
C9 4bitadder_1/fulladder_3/XOR_0/w_16_n1# 4bitadder_1/fulladder_3/XOR_0/bbar 0.03fF
C10 enable_0/and_5/a_n26_14# enable_0/and_5/w_26_9# 0.09fF
C11 comparator_0/4input_AND_1/w_68_n95# comparator_0/a2xnorb2 0.16fF
C12 enable_1/and_2/w_26_9# vdd 0.03fF
C13 a3out_2 b2out_2 0.30fF
C14 comparator_0/b3 a2out_2 0.48fF
C15 a2 b0 0.25fF
C16 comparator_0/3input_AND_1/not_0/in comparator_0/3input_AND_1/not_0/w_n2_10# 0.09fF
C17 4bitadder_0/fulladder_3/XOR_0/w_n34_n1# 4bitadder_0/fulladder_3/XOR_0/abar 0.03fF
C18 4bitadder_0/fulladder_3/XOR_0/w_16_n1# 4bitadder_0/fulladder_3/XOR_0/bbar 0.03fF
C19 enable_1/and_3/w_26_9# a3out_1 0.03fF
C20 comparator_0/4input_AND_2/not_0/in comparator_0/4input_AND_2/w_n8_2# 0.02fF
C21 b0 enable_2/and_4/w_n43_8# 0.09fF
C22 b1out_1 b3out_1 0.25fF
C23 decoder_0/and_3/w_n43_8# decoder_0/and_3/a_n26_14# 0.02fF
C24 comparator_0/not_2/w_n2_10# vdd 0.18fF
C25 enable_0/and_4/w_n43_8# b0 0.09fF
C26 b0 vdd 0.47fF
C27 vdd decoder_0/and_1/w_26_9# 0.03fF
C28 4bitadder_0/fulladder_0/and_1/w_26_9# vdd 0.03fF
C29 comparator_0/4input_AND_2/not_0/in comparator_0/a2xnorb2 0.18fF
C30 vdd s0 0.73fF
C31 comparator_0/4input_OR_0/w_n58_n43# vdd 0.03fF
C32 4bitadder_0/fulladder_0/or_0/w_58_101# 4bitadder_0/fulladder_0/or_0/a_n15_32# 0.13fF
C33 a3out_3 b0out_3 0.14fF
C34 comparator_0/a1bar comparator_0/a2xnorb2 0.26fF
C35 b2out_2 comparator_0/3input_AND_1/w_32_n21# 0.16fF
C36 4bitadder_0/fulladder_0/or_0/b gnd 0.37fF
C37 a3out_1 b2out_1 0.05fF
C38 vdd s0_sub 0.19fF
C39 4bitadder_1/fulladder_1/or_0/w_58_101# 4bitadder_1/fulladder_1/or_0/a_n15_32# 0.13fF
C40 4bitadder_0/fulladder_0/axorb vdd 0.15fF
C41 vdd 4bitadder_1/fulladder_2/XOR_1/w_n34_n1# 0.02fF
C42 4bitadder_0/fulladder_0/XOR_1/w_16_n1# s0 0.11fF
C43 enable_3/and_4/w_26_9# b0out_3 0.03fF
C44 a2out_2 a1out_2 0.75fF
C45 4bitadder_0/fulladder_0/and_0/w_26_9# vdd 0.03fF
C46 enable_0/and_7/a_n26_14# b3 0.31fF
C47 a0out_2 boout_2 0.87fF
C48 comparator_0/xnor_3/XOR_0/w_16_n1# comparator_0/xnor_3/XOR_0/bbar 0.03fF
C49 comparator_0/xnor_3/XOR_0/w_62_n20# comparator_0/xnor_3/not_0/in 0.04fF
C50 enable_1/en b0 0.28fF
C51 enable_1/en decoder_0/and_1/w_26_9# 0.03fF
C52 4bitadder_1/fulladder_0/and_1/w_n43_8# 4bitadder_1/b0xorM 0.09fF
C53 b0out_1 s0 0.17fF
C54 enable_2/a0 vdd 0.10fF
C55 a2out_1 4bitadder_1/fulladder_2/and_1/a_n26_14# 0.10fF
C56 4bitadder_1/fulladder_1/or_0/a_n15_32# 4bitadder_1/fulladder_1/or_0/b 0.19fF
C57 decoder_0/and_1/a_n26_14# decoder_0/and_1/b 0.29fF
C58 4bitadder_0/fulladder_0/XOR_1/abar s0 0.27fF
C59 4bitadder_0/fulladder_1/XOR_0/abar a1out_0 0.13fF
C60 4bitadder_1/fulladder_3/axorb 4bitadder_1/fulladder_3/XOR_1/w_62_37# 0.02fF
C61 4bitadder_1/c3 4bitadder_1/fulladder_3/XOR_1/w_16_n1# 0.11fF
C62 4bitadder_0/fulladder_3/or_0/a 4bitadder_0/fulladder_3/or_0/w_n48_101# 0.12fF
C63 gnd decoder_0/and_2/a 0.18fF
C64 4bitadder_0/fulladder_0/axorb 4bitadder_0/fulladder_0/XOR_1/abar 0.13fF
C65 comparator_0/5input_AND_1/not_0/in comparator_0/5input_AND_1/w_n4_n20# 0.03fF
C66 vdd 4bitadder_1/fulladder_3/and_0/w_n43_8# 0.07fF
C67 a0_out1 gnd 0.56fF
C68 4bitadder_1/fulladder_2/or_0/a_n15_32# 4bitadder_1/fulladder_2/or_0/b 0.19fF
C69 4bitadder_1/c3 4bitadder_1/fulladder_3/XOR_1/abar 0.27fF
C70 4bitadder_0/fulladder_1/XOR_0/w_16_n1# 4bitadder_0/fulladder_1/XOR_0/bbar 0.03fF
C71 enable_3/en a0 0.23fF
C72 4bitadder_0/fulladder_2/and_1/w_26_9# 4bitadder_0/fulladder_2/and_1/a_n26_14# 0.09fF
C73 4bitadder_1/fulladder_3/and_0/a_n26_14# 4bitadder_1/fulladder_3/and_0/w_n43_8# 0.02fF
C74 b0out_0 4bitadder_0/XOR_0/w_62_37# 0.02fF
C75 enable_1/and_7/w_n43_8# enable_1/and_7/a_n26_14# 0.02fF
C76 4bitadder_1/XOR_1/out s0 0.15fF
C77 4bitadder_0/fulladder_1/XOR_1/w_62_n20# 4bitadder_0/fulladder_1/XOR_1/abar 0.02fF
C78 b3out_1 4bitadder_1/XOR_3/abar 0.13fF
C79 4bitadder_1/c2 a2out_1 0.50fF
C80 vdd b1out_1 0.13fF
C81 comparator_0/a1xnorb1 comparator_0/5input_AND_1/w_31_n55# 0.21fF
C82 comparator_0/4input_OR_0/w_n58_n43# comparator_0/t6 0.13fF
C83 enable_3/and_7/a_n26_14# b3 0.31fF
C84 enable_3/and_5/a_n26_14# enable_3/and_5/w_26_9# 0.09fF
C85 b2 a1 0.31fF
C86 vdd 4bitadder_1/fulladder_1/and_0/w_n43_8# 0.07fF
C87 4bitadder_0/XOR_1/w_16_n1# vdd 0.02fF
C88 enable_2/and_3/w_n43_8# enable_2/and_3/a_n26_14# 0.02fF
C89 enable_0/and_2/a_n26_14# a2 0.31fF
C90 b3out_0 gnd 0.70fF
C91 4bitadder_0/XOR_2/abar gnd 0.13fF
C92 decoder_0/and_2/w_n43_8# decoder_0/and_2/a_n26_14# 0.02fF
C93 enable_1/and_1/w_n43_8# enable_1/and_1/a_n26_14# 0.02fF
C94 comparator_0/t8 comparator_0/t7 0.15fF
C95 4bitadder_0/XOR_0/abar gnd 0.15fF
C96 4bitadder_1/fulladder_1/XOR_1/w_62_n20# 4bitadder_1/fulladder_1/XOR_1/abar 0.02fF
C97 vdd comparator_0/4input_AND_0/w_68_n95# 0.02fF
C98 4bitadder_0/c2 a2out_0 0.50fF
C99 comparator_0/b2bar gnd 0.14fF
C100 comparator_0/3input_AND_1/not_0/in comparator_0/3input_AND_1/w_n14_24# 0.03fF
C101 enable_0/and_3/w_n43_8# enable_0/and_3/a_n26_14# 0.02fF
C102 AND_Block_0/and_3/w_n43_8# vdd 0.07fF
C103 4bitadder_1/fulladder_3/and_1/w_26_9# 4bitadder_1/fulladder_3/and_1/a_n26_14# 0.09fF
C104 comparator_0/4input_AND_0/w_n47_52# comparator_0/a3xnorb3 0.16fF
C105 gnd 4bitadder_1/fulladder_3/XOR_0/abar 0.15fF
C106 enable_1/and_4/w_26_9# vdd 0.03fF
C107 a0_out1 4bitadder_1/fulladder_0/XOR_0/w_62_37# 0.02fF
C108 comparator_0/xnor_1/XOR_0/w_62_37# b2out_2 0.13fF
C109 decoder_0/not_0/w_n2_10# decoder_0/and_2/a 0.03fF
C110 4bitadder_1/fulladder_1/XOR_0/bbar 4bitadder_1/fulladder_1/XOR_0/w_62_n20# 0.13fF
C111 comparator_0/3input_AND_1/not_0/in comparator_0/a3xnorb3 0.19fF
C112 4bitadder_0/fulladder_3/and_1/w_26_9# 4bitadder_0/fulladder_3/and_1/a_n26_14# 0.09fF
C113 4bitadder_1/XOR_3/out s0 0.16fF
C114 comparator_0/5input_AND_1/w_68_n82# comparator_0/a2xnorb2 0.16fF
C115 4bitadder_1/fulladder_0/and_1/w_n43_8# 4bitadder_1/fulladder_0/and_1/a_n26_14# 0.02fF
C116 vdd 4bitadder_1/fulladder_2/and_1/w_n43_8# 0.07fF
C117 4bitadder_1/fulladder_2/XOR_0/w_62_37# 4bitadder_1/XOR_2/out 0.13fF
C118 enable_0/and_7/w_26_9# b3out_0 0.03fF
C119 vdd a0out_2 0.68fF
C120 4bitadder_1/fulladder_0/and_0/a_n26_14# 4bitadder_1/fulladder_0/and_0/w_n43_8# 0.02fF
C121 b2out_2 comparator_0/xnor_1/not_0/in 0.13fF
C122 a2out_2 comparator_0/xnor_1/XOR_0/abar 0.13fF
C123 decoder_0/and_1/b decoder_0/and_1/w_n43_8# 0.09fF
C124 enable_1/and_4/w_26_9# b0out_1 0.03fF
C125 a0out_0 4bitadder_0/fulladder_0/and_1/a_n26_14# 0.10fF
C126 4bitadder_1/fulladder_1/axorb 4bitadder_1/fulladder_1/XOR_0/w_62_n20# 0.04fF
C127 s0_sub s0 0.04fF
C128 comparator_0/t1 gnd 0.01fF
C129 comparator_0/xnor_3/XOR_0/abar gnd 0.14fF
C130 4bitadder_0/fulladder_0/axorb s0 0.54fF
C131 comparator_0/a0xnorb0 comparator_0/4input_AND_0/not_0/in 0.18fF
C132 vdd 4bitadder_1/XOR_3/w_16_n1# 0.02fF
C133 enable_2/and_1/w_26_9# vdd 0.03fF
C134 comparator_0/t8 comparator_0/5input_AND_0/not_0/w_n2_10# 0.03fF
C135 4bitadder_1/fulladder_3/or_0/w_n48_101# 4bitadder_1/fulladder_3/or_0/a 0.12fF
C136 comparator_0/3input_AND_0/not_0/in comparator_0/3input_AND_0/w_32_n21# 0.02fF
C137 enable_2/and_0/w_26_9# vdd 0.03fF
C138 enable_0/en enable_0/and_6/w_n43_8# 0.09fF
C139 comparator_0/4input_AND_0/w_n8_2# comparator_0/a2xnorb2 0.16fF
C140 b2out_0 4bitadder_0/XOR_2/w_62_37# 0.02fF
C141 4bitadder_0/fulladder_2/or_0/a vdd 0.14fF
C142 decoder_0/and_1/b decoder_0/and_2/a 0.34fF
C143 comparator_0/xnor_3/XOR_0/w_62_37# a0out_2 0.02fF
C144 a1out_0 a2out_0 2.80fF
C145 comparator_0/4input_OR_1/w_n58_n43# comparator_0/t1 0.13fF
C146 comparator_0/a2xnorb2 comparator_0/b2bar 0.11fF
C147 b3 gnd 0.29fF
C148 gnd 4bitadder_1/c2 0.97fF
C149 comparator_0/xnor_0/XOR_0/w_n34_n1# a3out_2 0.11fF
C150 4bitadder_0/fulladder_2/or_0/a_n15_32# 4bitadder_0/fulladder_2/or_0/b 0.19fF
C151 vdd 4bitadder_1/fulladder_2/axorb 0.15fF
C152 4bitadder_1/fulladder_2/axorb 4bitadder_1/fulladder_2/XOR_0/w_62_n20# 0.04fF
C153 4bitadder_0/c2 vdd 0.17fF
C154 comparator_0/xnor_3/not_0/w_n2_10# comparator_0/xnor_3/not_0/in 0.09fF
C155 enable_3/and_2/w_26_9# a2out_3 0.03fF
C156 4bitadder_1/b0xorM 4bitadder_1/fulladder_0/XOR_0/bbar 0.02fF
C157 comparator_0/xnor_0/XOR_0/w_62_n20# comparator_0/xnor_0/XOR_0/abar 0.02fF
C158 enable_3/and_2/w_26_9# enable_3/and_2/a_n26_14# 0.09fF
C159 4bitadder_0/fulladder_2/or_0/a_n15_32# 4bitadder_0/fulladder_2/or_0/w_58_101# 0.13fF
C160 4bitadder_0/c1 4bitadder_0/fulladder_1/XOR_1/w_16_n1# 0.11fF
C161 b1out_1 s0 0.18fF
C162 4bitadder_0/fulladder_2/and_0/w_26_9# 4bitadder_0/fulladder_2/or_0/a 0.03fF
C163 4bitadder_0/XOR_1/w_16_n1# s0 0.11fF
C164 4bitadder_0/c1 4bitadder_0/fulladder_1/XOR_1/abar 0.27fF
C165 4bitadder_0/fulladder_0/or_0/a vdd 0.14fF
C166 4bitadder_1/fulladder_0/or_0/b 4bitadder_1/fulladder_0/or_0/w_n48_101# 0.12fF
C167 a3 enable_2/and_3/a_n26_14# 0.31fF
C168 b2 a3 0.31fF
C169 enable_1/and_3/w_n43_8# vdd 0.07fF
C170 s0_sub 4bitadder_1/fulladder_0/XOR_1/w_62_n20# 0.04fF
C171 b2out_2 comparator_0/3input_AND_1/not_0/in 0.19fF
C172 enable_2/and_4/w_n43_8# enable_2/and_4/a_n26_14# 0.02fF
C173 enable_0/and_3/a_n26_14# a3 0.31fF
C174 comparator_0/5input_AND_0/not_0/in gnd 0.10fF
C175 comparator_0/4input_OR_0/y comparator_0/t7 0.18fF
C176 comparator_0/5input_AND_0/not_0/in comparator_0/5input_AND_0/w_68_n82# 0.02fF
C177 vdd comparator_0/xnor_1/not_0/w_n2_10# 0.18fF
C178 4bitadder_0/fulladder_1/or_0/w_58_101# 4bitadder_0/c2 0.02fF
C179 vdd 4bitadder_1/fulladder_2/XOR_0/w_n34_n1# 0.02fF
C180 enable_3/en a1 0.25fF
C181 enable_1/and_0/a_n26_14# a0 0.31fF
C182 comparator_0/b3 a1out_2 0.82fF
C183 a3out_2 b1out_2 0.60fF
C184 vdd 4bitadder_1/fulladder_3/XOR_1/w_16_n1# 0.02fF
C185 enable_0/and_4/w_n43_8# enable_0/and_4/a_n26_14# 0.02fF
C186 AND_Block_0/and_2/a_n26_14# AND_Block_0/and_2/w_n43_8# 0.02fF
C187 b2 enable_3/and_6/w_n43_8# 0.09fF
C188 vdd comparator_0/3input_AND_1/w_69_n71# 0.03fF
C189 4bitadder_1/fulladder_2/XOR_0/w_62_n20# 4bitadder_1/fulladder_2/XOR_0/bbar 0.13fF
C190 enable_1/en enable_1/and_3/w_n43_8# 0.09fF
C191 4bitadder_1/fulladder_3/axorb 4bitadder_1/fulladder_3/XOR_0/w_62_37# 0.02fF
C192 gnd comparator_0/a3xnorb3 0.82fF
C193 vdd comparator_0/4input_AND_1/w_68_n95# 0.02fF
C194 enable_1/and_6/a_n26_14# enable_1/and_6/w_n43_8# 0.02fF
C195 a1out_0 vdd 0.28fF
C196 AND_Block_0/and_2/a_n26_14# AND_Block_0/and_2/w_26_9# 0.09fF
C197 s0_add vdd 0.19fF
C198 4bitadder_0/fulladder_3/or_0/w_58_101# fc_add 0.02fF
C199 b0out_3 gnd 0.22fF
C200 enable_3/and_0/w_n43_8# a0 0.09fF
C201 comparator_0/b0bar comparator_0/5input_AND_0/not_0/in 0.23fF
C202 4bitadder_0/fulladder_1/and_1/w_n43_8# 4bitadder_0/XOR_1/out 0.09fF
C203 enable_0/en enable_0/and_0/w_n43_8# 0.09fF
C204 s0 4bitadder_1/XOR_3/w_16_n1# 0.11fF
C205 vdd 4bitadder_1/XOR_0/w_n34_n1# 0.02fF
C206 vdd 4bitadder_1/fulladder_0/XOR_1/w_n34_n1# 0.02fF
C207 comparator_0/a1xnorb1 gnd 1.03fF
C208 4bitadder_0/fulladder_3/axorb vdd 0.15fF
C209 enable_1/and_6/a_n26_14# enable_1/and_6/w_26_9# 0.09fF
C210 4bitadder_0/fulladder_1/or_0/a gnd 0.01fF
C211 decoder_0/and_0/w_n43_8# decoder_0/and_1/b 0.09fF
C212 comparator_0/xnor_2/XOR_0/w_16_n1# b1out_2 0.11fF
C213 4bitadder_0/fulladder_0/or_0/w_58_101# 4bitadder_0/c1 0.02fF
C214 out0 gnd 0.01fF
C215 comparator_0/4input_AND_0/not_0/w_n2_10# comparator_0/4input_AND_0/not_0/in 0.09fF
C216 s0 4bitadder_1/XOR_3/abar 0.30fF
C217 gnd 4bitadder_1/fulladder_0/or_0/a 0.01fF
C218 AND_Block_0/and_0/w_26_9# vdd 0.03fF
C219 4bitadder_0/c1 gnd 0.77fF
C220 vdd comparator_0/a1bar 0.22fF
C221 4bitadder_0/fulladder_2/or_0/a_n15_32# 4bitadder_0/fulladder_2/or_0/w_n48_101# 0.05fF
C222 a1out_1 b2out_1 0.25fF
C223 b0out_1 4bitadder_1/XOR_0/w_n34_n1# 0.11fF
C224 enable_1/and_5/w_26_9# vdd 0.03fF
C225 comparator_0/b0bar comparator_0/a3xnorb3 0.28fF
C226 b1out_2 comparator_0/xnor_2/XOR_0/abar 0.30fF
C227 enable_2/and_7/w_n43_8# enable_2/and_7/a_n26_14# 0.02fF
C228 enable_3/and_0/w_26_9# a0out_3 0.03fF
C229 comparator_0/t4 comparator_0/t3 0.19fF
C230 comparator_0/4input_AND_0/not_0/in comparator_0/4input_AND_0/w_29_n46# 0.02fF
C231 comparator_0/5input_AND_0/not_0/in comparator_0/a2xnorb2 0.23fF
C232 4bitadder_1/fulladder_0/and_0/w_26_9# 4bitadder_1/fulladder_0/or_0/a 0.03fF
C233 4bitadder_0/fulladder_1/XOR_0/w_62_37# 4bitadder_0/XOR_1/out 0.13fF
C234 vdd 4bitadder_1/fulladder_2/or_0/w_n48_101# 0.05fF
C235 comparator_0/b0bar comparator_0/a1xnorb1 0.29fF
C236 comparator_0/4input_OR_1/y comparator_0/t3 0.18fF
C237 a2out_3 a3out_3 0.39fF
C238 a1out_1 4bitadder_1/fulladder_1/and_1/a_n26_14# 0.10fF
C239 4bitadder_0/c3 4bitadder_0/XOR_3/out 0.41fF
C240 4bitadder_1/fulladder_2/axorb 4bitadder_1/fulladder_2/XOR_1/w_n34_n1# 0.11fF
C241 enable_1/and_0/w_n43_8# vdd 0.07fF
C242 enable_0/and_6/w_n43_8# vdd 0.07fF
C243 a3 enable_2/a2 0.10fF
C244 4bitadder_0/XOR_3/w_n34_n1# vdd 0.02fF
C245 a3out_2 a2out_2 0.63fF
C246 comparator_0/a2xnorb2 comparator_0/a3xnorb3 7.69fF
C247 enable_3/and_3/w_26_9# enable_3/and_3/a_n26_14# 0.09fF
C248 decoder_0/and_2/w_n43_8# s1 0.09fF
C249 4bitadder_1/XOR_1/out 4bitadder_1/fulladder_1/XOR_0/abar 0.25fF
C250 4bitadder_1/fulladder_0/XOR_0/w_n34_n1# a0_out1 0.11fF
C251 enable_1/and_7/w_n43_8# b3 0.09fF
C252 4bitadder_0/fulladder_1/axorb 4bitadder_0/c1 0.54fF
C253 4bitadder_0/fulladder_3/and_0/a_n26_14# 4bitadder_0/fulladder_3/and_0/w_26_9# 0.09fF
C254 vdd 4bitadder_1/fulladder_3/and_1/w_26_9# 0.03fF
C255 comparator_0/a1xnorb1 comparator_0/a2xnorb2 1.39fF
C256 4bitadder_0/XOR_2/out 4bitadder_0/XOR_2/w_62_n20# 0.04fF
C257 enable_1/and_0/w_n43_8# enable_1/en 0.09fF
C258 a3out_0 a0_out1 0.21fF
C259 comparator_0/t7 comparator_0/4input_AND_1/not_0/w_n2_10# 0.03fF
C260 vdd comparator_0/xnor_1/XOR_0/w_n34_n1# 0.02fF
C261 4bitadder_0/fulladder_0/XOR_0/w_62_n20# 4bitadder_0/fulladder_0/XOR_0/bbar 0.13fF
C262 enable_2/and_1/w_n43_8# vdd 0.07fF
C263 4bitadder_0/fulladder_0/or_0/a 4bitadder_0/fulladder_0/and_0/w_26_9# 0.03fF
C264 b0 enable_2/and_4/a_n26_14# 0.31fF
C265 gnd 4bitadder_1/fulladder_3/or_0/b 0.37fF
C266 b2out_2 gnd 0.98fF
C267 enable_0/and_4/a_n26_14# b0 0.31fF
C268 a0out_0 gnd 0.46fF
C269 vdd decoder_0/and_1/w_n43_8# 0.07fF
C270 enable_2/and_6/w_n43_8# vdd 0.07fF
C271 gnd 4bitadder_1/XOR_1/abar 0.23fF
C272 comparator_0/4input_AND_2/w_29_n46# comparator_0/a2xnorb2 0.16fF
C273 a3out_2 comparator_0/not_7/w_n2_10# 0.09fF
C274 4bitadder_0/fulladder_0/XOR_1/w_62_37# s0 0.13fF
C275 enable_3/en a3 0.23fF
C276 enable_0/en b3 0.10fF
C277 enable_2/en gnd 0.16fF
C278 comparator_0/xnor_3/XOR_0/w_16_n1# boout_2 0.11fF
C279 4bitadder_0/fulladder_0/axorb 4bitadder_0/fulladder_0/XOR_1/w_62_37# 0.02fF
C280 enable_3/and_1/w_n43_8# enable_3/en 0.09fF
C281 a1out_0 s0 2.21fF
C282 enable_2/and_6/w_26_9# vdd 0.03fF
C283 b3out_0 a3out_0 0.11fF
C284 decoder_0/and_1/a_n26_14# decoder_0/and_1/w_26_9# 0.09fF
C285 4bitadder_1/XOR_2/out a2out_1 1.88fF
C286 4bitadder_1/fulladder_2/and_1/w_26_9# 4bitadder_1/fulladder_2/or_0/b 0.03fF
C287 s0_add s0 0.04fF
C288 4bitadder_1/c3 4bitadder_1/fulladder_3/XOR_1/w_62_37# 0.13fF
C289 4bitadder_0/fulladder_2/XOR_1/w_n34_n1# vdd 0.02fF
C290 4bitadder_0/fulladder_1/XOR_0/bbar 4bitadder_0/XOR_1/out 0.02fF
C291 enable_3/and_7/w_26_9# vdd 0.03fF
C292 enable_2/and_7/w_26_9# enable_2/and_7/a_n26_14# 0.09fF
C293 enable_3/and_6/w_n43_8# enable_3/en 0.09fF
C294 enable_3/and_5/w_n43_8# enable_3/and_5/a_n26_14# 0.02fF
C295 boout_2 comparator_0/xnor_3/XOR_0/abar 0.30fF
C296 vdd decoder_0/and_2/a 0.04fF
C297 vdd comparator_0/5input_AND_1/w_68_n82# 0.05fF
C298 4bitadder_1/XOR_3/w_62_37# b3out_1 0.02fF
C299 4bitadder_1/c3 s3_sub 0.04fF
C300 vdd a0_out1 0.26fF
C301 a2out_2 comparator_0/b3bar 0.21fF
C302 enable_2/and_0/w_26_9# a0out_2 0.03fF
C303 enable_3/and_5/a_n26_14# b1 0.31fF
C304 4bitadder_0/fulladder_2/and_1/w_n43_8# a2out_0 0.09fF
C305 vdd 4bitadder_1/fulladder_1/XOR_0/w_16_n1# 0.02fF
C306 4bitadder_0/fulladder_1/and_0/w_26_9# 4bitadder_0/fulladder_1/or_0/a 0.03fF
C307 s0 s1 1.27fF
C308 4bitadder_0/fulladder_3/XOR_1/w_n34_n1# vdd 0.02fF
C309 4bitadder_0/fulladder_1/XOR_1/w_n34_n1# 4bitadder_0/fulladder_1/XOR_1/abar 0.03fF
C310 4bitadder_0/fulladder_1/XOR_1/w_16_n1# 4bitadder_0/fulladder_1/XOR_1/bbar 0.03fF
C311 4bitadder_0/fulladder_1/XOR_1/w_62_n20# s1_add 0.04fF
C312 4bitadder_1/XOR_3/w_62_n20# 4bitadder_1/XOR_3/bbar 0.13fF
C313 enable_0/and_0/w_n43_8# vdd 0.07fF
C314 4bitadder_0/XOR_2/w_16_n1# vdd 0.02fF
C315 4bitadder_1/fulladder_1/and_1/w_26_9# 4bitadder_1/fulladder_1/and_1/a_n26_14# 0.09fF
C316 vdd comparator_0/and_0/w_n43_8# 0.07fF
C317 4bitadder_0/XOR_3/w_62_n20# 4bitadder_0/XOR_3/bbar 0.13fF
C318 b3out_0 vdd 0.13fF
C319 b1 b3 0.24fF
C320 decoder_0/and_2/w_n43_8# decoder_0/and_2/a 0.09fF
C321 4bitadder_1/fulladder_1/XOR_1/w_n34_n1# 4bitadder_1/fulladder_1/XOR_1/abar 0.03fF
C322 4bitadder_1/fulladder_1/XOR_1/w_16_n1# 4bitadder_1/fulladder_1/XOR_1/bbar 0.03fF
C323 4bitadder_1/fulladder_1/XOR_1/w_62_n20# s1_sub 0.04fF
C324 vdd comparator_0/4input_AND_0/w_n8_2# 0.02fF
C325 4bitadder_0/fulladder_2/axorb 4bitadder_0/XOR_2/out 0.13fF
C326 4bitadder_0/fulladder_2/XOR_0/w_62_37# a2out_0 0.02fF
C327 vdd 4bitadder_1/fulladder_3/XOR_0/w_16_n1# 0.02fF
C328 b2out_3 AND_Block_0/and_2/a_n26_14# 0.31fF
C329 vdd comparator_0/b2bar 1.10fF
C330 enable_3/and_3/w_26_9# vdd 0.03fF
C331 4bitadder_1/fulladder_3/and_1/w_n43_8# a3out_1 0.09fF
C332 4bitadder_1/fulladder_0/and_0/a_n26_14# 4bitadder_1/fulladder_0/and_0/w_26_9# 0.09fF
C333 b2 enable_2/and_6/a_n26_14# 0.31fF
C334 decoder_0/and_2/a_n26_14# s1 0.31fF
C335 4bitadder_1/fulladder_2/or_0/a_n15_32# 4bitadder_1/fulladder_2/or_0/w_58_101# 0.13fF
C336 b0out_0 4bitadder_0/XOR_0/w_n34_n1# 0.11fF
C337 comparator_0/xnor_1/XOR_0/w_62_37# a2out_2 0.02fF
C338 4bitadder_0/XOR_3/bbar s0 0.02fF
C339 4bitadder_0/fulladder_3/and_1/w_n43_8# a3out_0 0.09fF
C340 enable_3/and_4/w_26_9# enable_3/and_4/a_n26_14# 0.09fF
C341 comparator_0/t4 comparator_0/t2 0.19fF
C342 comparator_0/4input_AND_1/not_0/in comparator_0/4input_AND_1/w_29_n46# 0.02fF
C343 4bitadder_0/fulladder_3/or_0/a gnd 0.01fF
C344 vdd 4bitadder_1/fulladder_1/XOR_0/w_n34_n1# 0.02fF
C345 vdd comparator_0/3input_AND_1/not_0/w_n2_10# 0.18fF
C346 4bitadder_1/fulladder_0/or_0/a_n15_32# 4bitadder_1/fulladder_0/or_0/w_n48_101# 0.05fF
C347 enable_0/and_7/w_n43_8# enable_0/and_7/a_n26_14# 0.02fF
C348 4bitadder_1/fulladder_1/XOR_0/w_16_n1# 4bitadder_1/XOR_1/out 0.11fF
C349 vdd comparator_0/xnor_3/XOR_0/w_16_n1# 0.02fF
C350 comparator_0/4input_OR_1/y comparator_0/t2 0.18fF
C351 comparator_0/xnor_1/XOR_0/w_62_n20# comparator_0/xnor_1/XOR_0/bbar 0.13fF
C352 gnd 4bitadder_1/XOR_2/out 0.42fF
C353 4bitadder_0/b0xorM a0out_0 1.79fF
C354 4bitadder_0/fulladder_0/and_1/w_26_9# 4bitadder_0/fulladder_0/or_0/b 0.03fF
C355 enable_1/and_5/w_26_9# b1out_1 0.03fF
C356 b2 enable_2/b1 0.11fF
C357 s0 decoder_0/and_1/w_n43_8# 0.09fF
C358 comparator_0/xnor_3/not_0/in gnd 0.03fF
C359 4bitadder_1/XOR_2/out 4bitadder_1/XOR_2/w_62_37# 0.02fF
C360 4bitadder_0/fulladder_2/and_1/w_n43_8# vdd 0.07fF
C361 4bitadder_1/fulladder_1/and_0/a_n26_14# 4bitadder_1/c1 0.10fF
C362 4bitadder_0/fulladder_1/and_0/w_n43_8# 4bitadder_0/fulladder_1/and_0/a_n26_14# 0.02fF
C363 a0 gnd 0.21fF
C364 b3 a2 0.21fF
C365 comparator_0/t3 comparator_0/t2 0.19fF
C366 boout_2 comparator_0/a3xnorb3 0.48fF
C367 vdd decoder_0/and_0/w_n43_8# 0.07fF
C368 vdd comparator_0/not_5/w_n2_10# 0.18fF
C369 enable_0/and_0/w_n43_8# enable_0/and_0/a_n26_14# 0.02fF
C370 enable_2/and_5/w_n43_8# enable_2/b1 0.09fF
C371 decoder_0/and_0/a_n26_14# decoder_0/and_0/w_26_9# 0.09fF
C372 4bitadder_1/fulladder_2/XOR_1/w_62_37# s2_sub 0.02fF
C373 4bitadder_1/b0xorM gnd 0.42fF
C374 comparator_0/a1xnorb1 boout_2 0.85fF
C375 enable_1/and_5/w_n43_8# b1 0.09fF
C376 s0 decoder_0/and_2/a 0.12fF
C377 4bitadder_0/fulladder_3/and_1/w_n43_8# vdd 0.07fF
C378 4bitadder_0/fulladder_0/and_0/a_n26_14# 4bitadder_0/fulladder_0/and_0/w_n43_8# 0.02fF
C379 b3 vdd 0.34fF
C380 vdd 4bitadder_1/c2 0.17fF
C381 a0_out1 s0 0.29fF
C382 comparator_0/not_0/w_n2_10# comparator_0/b0bar 0.03fF
C383 comparator_0/and_1/w_26_9# comparator_0/and_1/a_n26_14# 0.09fF
C384 4bitadder_0/fulladder_2/XOR_0/abar 4bitadder_0/XOR_2/out 0.25fF
C385 comparator_0/b1bar gnd 0.14fF
C386 a3out_2 comparator_0/b3 3.20fF
C387 comparator_0/xnor_0/XOR_0/w_n34_n1# comparator_0/xnor_0/XOR_0/abar 0.03fF
C388 comparator_0/xnor_0/XOR_0/w_16_n1# comparator_0/xnor_0/XOR_0/bbar 0.03fF
C389 comparator_0/xnor_0/XOR_0/w_62_n20# comparator_0/xnor_0/not_0/in 0.04fF
C390 enable_3/and_2/w_n43_8# a2 0.09fF
C391 4bitadder_1/c1 4bitadder_1/fulladder_1/XOR_1/w_16_n1# 0.11fF
C392 4bitadder_0/fulladder_1/axorb 4bitadder_0/fulladder_1/XOR_1/w_n34_n1# 0.11fF
C393 4bitadder_0/c1 4bitadder_0/fulladder_1/XOR_1/w_62_37# 0.13fF
C394 4bitadder_1/fulladder_1/or_0/w_58_101# 4bitadder_1/c2 0.02fF
C395 4bitadder_0/XOR_2/w_16_n1# s0 0.11fF
C396 4bitadder_0/c3 4bitadder_0/fulladder_3/XOR_1/w_16_n1# 0.11fF
C397 enable_1/en b3 0.21fF
C398 b2 enable_2/a2 0.10fF
C399 4bitadder_1/fulladder_2/and_0/a_n26_14# 4bitadder_1/c2 0.10fF
C400 4bitadder_1/c1 4bitadder_1/fulladder_1/XOR_1/abar 0.27fF
C401 4bitadder_0/c1 s1_add 0.04fF
C402 enable_3/and_2/w_n43_8# vdd 0.07fF
C403 4bitadder_1/fulladder_3/XOR_0/w_n34_n1# a3out_1 0.11fF
C404 4bitadder_1/fulladder_3/XOR_0/w_16_n1# 4bitadder_1/XOR_3/out 0.11fF
C405 comparator_0/not_2/w_n2_10# comparator_0/b2bar 0.03fF
C406 4bitadder_0/fulladder_2/XOR_1/w_62_n20# 4bitadder_0/fulladder_2/XOR_1/bbar 0.13fF
C407 b3out_0 s0 0.51fF
C408 a2out_3 gnd 0.17fF
C409 gnd 4bitadder_1/fulladder_3/or_0/a 0.01fF
C410 4bitadder_0/fulladder_1/or_0/w_n48_101# 4bitadder_0/fulladder_1/or_0/a_n15_32# 0.05fF
C411 enable_3/and_7/w_n43_8# b3 0.09fF
C412 4bitadder_0/XOR_2/abar s0 0.28fF
C413 4bitadder_0/c3 4bitadder_0/fulladder_3/XOR_1/abar 0.27fF
C414 4bitadder_0/fulladder_3/XOR_0/w_n34_n1# a3out_0 0.11fF
C415 4bitadder_0/fulladder_3/XOR_0/w_16_n1# 4bitadder_0/XOR_3/out 0.11fF
C416 a2out_3 AND_Block_0/and_2/w_n43_8# 0.09fF
C417 4bitadder_0/XOR_0/abar s0 1.07fF
C418 comparator_0/5input_AND_0/not_0/in comparator_0/5input_AND_0/w_n4_n20# 0.03fF
C419 4bitadder_1/fulladder_3/XOR_0/abar 4bitadder_1/XOR_3/out 0.25fF
C420 4bitadder_1/fulladder_0/axorb 4bitadder_1/fulladder_0/and_0/w_n43_8# 0.09fF
C421 enable_2/en enable_2/and_2/w_n43_8# 0.09fF
C422 a3out_2 a1out_2 0.75fF
C423 4bitadder_1/b0xorM 4bitadder_1/fulladder_0/XOR_0/w_62_37# 0.13fF
C424 4bitadder_0/fulladder_3/XOR_0/abar 4bitadder_0/XOR_3/out 0.25fF
C425 vdd comparator_0/3input_AND_1/w_n14_24# 0.03fF
C426 vdd comparator_0/5input_AND_0/w_106_n113# 0.04fF
C427 AND_Block_0/and_3/a_n26_14# b3out_3 0.31fF
C428 vdd 4bitadder_1/XOR_2/w_n34_n1# 0.02fF
C429 AND_Block_0/and_0/w_n43_8# vdd 0.07fF
C430 a2out_1 a3out_1 11.02fF
C431 vdd comparator_0/4input_AND_1/w_n8_2# 0.02fF
C432 vdd s3_sub 0.10fF
C433 comparator_0/3input_AND_1/w_n14_24# comparator_0/a2bar 0.16fF
C434 vdd comparator_0/xnor_2/XOR_0/w_n34_n1# 0.02fF
C435 b2 enable_3/en 0.23fF
C436 4bitadder_1/XOR_3/out 4bitadder_1/XOR_3/w_62_37# 0.02fF
C437 4bitadder_1/fulladder_0/XOR_1/w_16_n1# vdd 0.02fF
C438 4bitadder_1/fulladder_3/XOR_1/w_62_n20# 4bitadder_1/fulladder_3/XOR_1/bbar 0.13fF
C439 vdd comparator_0/a3xnorb3 1.70fF
C440 enable_1/and_5/w_n43_8# vdd 0.07fF
C441 vdd decoder_0/and_2/w_26_9# 0.03fF
C442 b2out_2 boout_2 0.30fF
C443 comparator_0/b1bar comparator_0/a2xnorb2 0.51fF
C444 b0out_3 vdd 0.16fF
C445 4bitadder_0/XOR_3/out 4bitadder_0/XOR_3/w_62_37# 0.02fF
C446 b1out_2 gnd 1.06fF
C447 s0 4bitadder_1/XOR_3/w_62_37# 0.13fF
C448 gnd 4bitadder_1/fulladder_1/or_0/a 0.01fF
C449 4bitadder_0/fulladder_3/XOR_1/w_62_n20# 4bitadder_0/fulladder_3/XOR_1/bbar 0.13fF
C450 comparator_0/a2bar comparator_0/a3xnorb3 0.19fF
C451 4bitadder_0/fulladder_0/XOR_1/w_62_37# s0_add 0.02fF
C452 4bitadder_1/c1 gnd 0.77fF
C453 vdd 4bitadder_1/fulladder_1/and_1/w_n43_8# 0.07fF
C454 vdd comparator_0/a1xnorb1 0.87fF
C455 comparator_0/xnor_2/XOR_0/w_62_37# b1out_2 0.13fF
C456 4bitadder_0/fulladder_1/or_0/a vdd 0.14fF
C457 vdd comparator_0/not_1/w_n2_10# 0.18fF
C458 4bitadder_0/fulladder_3/XOR_0/w_n34_n1# vdd 0.02fF
C459 vdd comparator_0/4input_AND_2/not_0/w_n2_10# 0.18fF
C460 a1out_3 b0out_3 0.21fF
C461 b2out_1 4bitadder_1/XOR_2/abar 0.13fF
C462 4bitadder_1/XOR_0/bbar 4bitadder_1/XOR_0/w_16_n1# 0.03fF
C463 enable_1/and_5/w_n43_8# enable_1/en 0.09fF
C464 vdd 4bitadder_1/fulladder_0/or_0/a 0.14fF
C465 4bitadder_1/fulladder_0/XOR_0/abar gnd 0.15fF
C466 comparator_0/t8 comparator_0/t5 0.21fF
C467 b1out_2 comparator_0/xnor_2/not_0/in 0.13fF
C468 a1out_2 comparator_0/xnor_2/XOR_0/abar 0.13fF
C469 4bitadder_0/c1 vdd 0.12fF
C470 b3 b0 0.35fF
C471 b1 enable_2/en 0.10fF
C472 comparator_0/4input_AND_0/not_0/in comparator_0/4input_AND_0/w_n47_52# 0.02fF
C473 boout_2 comparator_0/5input_AND_1/w_n4_n20# 0.18fF
C474 4bitadder_0/fulladder_3/or_0/a 4bitadder_0/fulladder_3/and_0/w_26_9# 0.03fF
C475 vdd comparator_0/4input_AND_2/w_29_n46# 0.02fF
C476 4bitadder_0/fulladder_1/XOR_0/w_16_n1# 4bitadder_0/XOR_1/out 0.11fF
C477 vdd 4bitadder_1/fulladder_0/XOR_0/w_16_n1# 0.02fF
C478 comparator_0/a3bar comparator_0/and_1/w_n43_8# 0.09fF
C479 4bitadder_0/XOR_0/bbar 4bitadder_0/XOR_0/w_16_n1# 0.03fF
C480 4bitadder_0/fulladder_3/axorb 4bitadder_0/fulladder_3/XOR_0/w_62_n20# 0.04fF
C481 enable_0/and_0/w_26_9# vdd 0.03fF
C482 4bitadder_1/c1 4bitadder_1/fulladder_0/or_0/w_58_101# 0.02fF
C483 b1out_2 comparator_0/4input_AND_2/w_n8_2# 0.16fF
C484 a1 gnd 0.27fF
C485 enable_2/and_0/a_n26_14# enable_2/and_0/w_n43_8# 0.02fF
C486 enable_3/and_3/w_n43_8# a3 0.09fF
C487 enable_1/and_1/w_n43_8# a1 0.09fF
C488 4bitadder_1/c2 4bitadder_1/fulladder_2/XOR_1/bbar 0.02fF
C489 4bitadder_1/XOR_1/out 4bitadder_1/fulladder_1/and_1/w_n43_8# 0.09fF
C490 4bitadder_0/fulladder_1/XOR_0/w_62_37# 4bitadder_0/fulladder_1/axorb 0.02fF
C491 b1out_2 comparator_0/a2xnorb2 0.26fF
C492 comparator_0/4input_AND_1/not_0/in comparator_0/4input_AND_1/not_0/w_n2_10# 0.09fF
C493 comparator_0/a0xnorb0 comparator_0/xnor_3/not_0/w_n2_10# 0.03fF
C494 enable_3/and_4/w_n43_8# vdd 0.07fF
C495 out1 gnd 0.01fF
C496 enable_0/en a0 0.38fF
C497 4bitadder_0/c2 4bitadder_0/fulladder_2/XOR_1/bbar 0.02fF
C498 4bitadder_0/fulladder_2/axorb 4bitadder_0/fulladder_2/XOR_1/abar 0.13fF
C499 gnd a3out_1 1.05fF
C500 a2out_2 gnd 0.88fF
C501 a2 enable_2/en 0.15fF
C502 4bitadder_1/fulladder_1/axorb 4bitadder_1/fulladder_1/XOR_0/w_62_37# 0.02fF
C503 b1out_0 4bitadder_0/XOR_1/abar 0.13fF
C504 enable_3/and_1/w_26_9# enable_3/and_1/a_n26_14# 0.09fF
C505 vdd b2out_2 1.44fF
C506 a0out_0 vdd 0.26fF
C507 enable_2/en enable_2/and_4/w_n43_8# 0.09fF
C508 4bitadder_0/fulladder_0/or_0/w_n48_101# vdd 0.05fF
C509 enable_0/and_2/w_26_9# a2out_0 0.03fF
C510 b2out_2 comparator_0/a2bar 0.27fF
C511 comparator_0/a0bar comparator_0/not_4/w_n2_10# 0.03fF
C512 4bitadder_0/fulladder_2/and_0/w_n43_8# vdd 0.07fF
C513 AND_Block_0/and_3/a_n26_14# AND_Block_0/and_3/w_26_9# 0.09fF
C514 4bitadder_1/fulladder_0/XOR_1/w_16_n1# s0 0.11fF
C515 enable_2/en vdd 1.03fF
C516 vdd 4bitadder_1/fulladder_3/and_0/w_26_9# 0.03fF
C517 4bitadder_1/fulladder_2/and_1/w_n43_8# 4bitadder_1/fulladder_2/and_1/a_n26_14# 0.02fF
C518 4bitadder_1/fulladder_0/XOR_1/w_62_37# s0 0.13fF
C519 4bitadder_0/fulladder_0/XOR_0/w_62_37# 4bitadder_0/b0xorM 0.13fF
C520 4bitadder_1/fulladder_1/and_0/w_26_9# 4bitadder_1/fulladder_1/or_0/a 0.03fF
C521 s0_sub 4bitadder_1/fulladder_0/XOR_1/w_62_37# 0.02fF
C522 a3out_3 b1out_3 0.11fF
C523 s0 4bitadder_1/XOR_2/bbar 0.02fF
C524 boout_2 comparator_0/xnor_3/not_0/in 0.13fF
C525 a0out_2 comparator_0/xnor_3/XOR_0/abar 0.13fF
C526 comparator_0/not_0/w_n2_10# boout_2 0.09fF
C527 4bitadder_0/fulladder_1/XOR_0/w_62_n20# 4bitadder_0/fulladder_1/XOR_0/bbar 0.13fF
C528 gnd 4bitadder_1/fulladder_2/XOR_1/abar 0.15fF
C529 AND_Block_0/and_1/w_n43_8# vdd 0.07fF
C530 decoder_0/and_1/a_n26_14# decoder_0/and_1/w_n43_8# 0.02fF
C531 4bitadder_1/fulladder_3/and_0/a_n26_14# 4bitadder_1/fulladder_3/and_0/w_26_9# 0.09fF
C532 vdd comparator_0/5input_AND_1/w_n4_n20# 0.05fF
C533 b1out_0 gnd 0.52fF
C534 enable_0/en enable_0/and_1/w_n43_8# 0.09fF
C535 enable_0/and_0/w_26_9# enable_0/and_0/a_n26_14# 0.09fF
C536 comparator_0/5input_AND_1/not_0/in comparator_0/5input_AND_1/w_106_n113# 0.03fF
C537 4bitadder_0/fulladder_1/XOR_0/w_n34_n1# 4bitadder_0/fulladder_1/XOR_0/abar 0.03fF
C538 comparator_0/4input_OR_0/y comparator_0/t5 0.18fF
C539 AND_Block_0/and_1/w_n43_8# a1out_3 0.09fF
C540 enable_0/and_6/w_26_9# b2out_0 0.03fF
C541 4bitadder_1/XOR_0/w_62_37# b0out_1 0.02fF
C542 a1 enable_3/and_1/a_n26_14# 0.31fF
C543 b1 a0 0.28fF
C544 4bitadder_1/fulladder_1/axorb 4bitadder_1/fulladder_1/XOR_1/abar 0.13fF
C545 a2out_0 4bitadder_0/fulladder_2/and_1/a_n26_14# 0.10fF
C546 decoder_0/and_2/w_26_9# decoder_0/and_2/a_n26_14# 0.09fF
C547 enable_1/and_1/w_26_9# a1out_1 0.03fF
C548 a2out_2 comparator_0/a2xnorb2 0.17fF
C549 a2out_3 b2out_3 2.92fF
C550 enable_1/and_2/w_n43_8# enable_1/and_2/a_n26_14# 0.02fF
C551 enable_0/en enable_0/and_5/w_n43_8# 0.09fF
C552 comparator_0/4input_AND_0/not_0/in gnd 0.03fF
C553 enable_2/and_2/w_26_9# vdd 0.03fF
C554 b3out_2 comparator_0/b3 0.10fF
C555 4bitadder_0/fulladder_2/XOR_0/w_62_n20# 4bitadder_0/fulladder_2/axorb 0.04fF
C556 vdd comparator_0/3input_AND_0/w_69_n71# 0.03fF
C557 b1out_0 4bitadder_0/XOR_1/w_62_37# 0.02fF
C558 4bitadder_0/fulladder_3/axorb 4bitadder_0/fulladder_3/XOR_1/w_n34_n1# 0.11fF
C559 enable_0/and_2/w_26_9# vdd 0.03fF
C560 comparator_0/4input_AND_1/not_0/in gnd 0.21fF
C561 decoder_0/and_2/a s1 0.24fF
C562 vdd comparator_0/t7 0.04fF
C563 4bitadder_0/XOR_0/w_16_n1# vdd 0.02fF
C564 enable_3/and_4/w_n43_8# b0 0.09fF
C565 a3 gnd 0.27fF
C566 comparator_0/4input_AND_1/not_0/in comparator_0/4input_AND_1/w_n47_52# 0.02fF
C567 a3out_1 4bitadder_1/fulladder_3/and_1/a_n26_14# 0.10fF
C568 comparator_0/not_2/w_n2_10# b2out_2 0.09fF
C569 4bitadder_0/fulladder_3/or_0/a vdd 0.14fF
C570 comparator_0/b3 comparator_0/and_1/a_n26_14# 0.10fF
C571 enable_0/and_7/w_n43_8# enable_0/en 0.09fF
C572 4bitadder_0/c3 4bitadder_0/fulladder_3/and_0/w_n43_8# 0.09fF
C573 4bitadder_1/c2 4bitadder_1/fulladder_2/axorb 0.54fF
C574 a3out_0 4bitadder_0/fulladder_3/and_1/a_n26_14# 0.10fF
C575 enable_2/and_4/w_26_9# boout_2 0.03fF
C576 4bitadder_0/fulladder_0/and_1/w_n43_8# 4bitadder_0/fulladder_0/and_1/a_n26_14# 0.02fF
C577 4bitadder_1/fulladder_1/axorb gnd 0.09fF
C578 a0 a2 0.40fF
C579 a0out_0 s0 0.55fF
C580 comparator_0/and_0/w_n43_8# comparator_0/and_0/a_n26_14# 0.02fF
C581 comparator_0/and_0/w_26_9# comparator_0/t5 0.03fF
C582 comparator_0/not_0/w_n2_10# vdd 0.18fF
C583 AND_Block_0/and_1/w_26_9# vdd 0.03fF
C584 s0 4bitadder_1/XOR_1/abar 0.25fF
C585 4bitadder_0/fulladder_1/XOR_1/w_n34_n1# vdd 0.02fF
C586 b0 enable_2/en 0.31fF
C587 4bitadder_1/fulladder_2/XOR_0/abar a2out_1 0.13fF
C588 a1out_1 4bitadder_1/fulladder_1/XOR_0/w_62_37# 0.02fF
C589 a0out_2 comparator_0/a3xnorb3 0.28fF
C590 4bitadder_0/XOR_2/out gnd 0.42fF
C591 4bitadder_0/fulladder_0/or_0/a_n15_32# 4bitadder_0/fulladder_0/or_0/b 0.19fF
C592 a2out_1 b2out_1 0.16fF
C593 a0 vdd 0.31fF
C594 4bitadder_1/c3 a3out_1 0.40fF
C595 vdd 4bitadder_1/fulladder_1/XOR_1/w_n34_n1# 0.02fF
C596 4bitadder_1/fulladder_1/XOR_0/w_n34_n1# 4bitadder_1/fulladder_1/XOR_0/abar 0.03fF
C597 b1 enable_0/and_5/w_n43_8# 0.09fF
C598 comparator_0/4input_AND_0/not_0/in comparator_0/a2xnorb2 0.18fF
C599 b1out_2 boout_2 0.73fF
C600 vdd comparator_0/5input_AND_0/not_0/w_n2_10# 0.17fF
C601 comparator_0/a1xnorb1 a0out_2 0.40fF
C602 4bitadder_1/XOR_0/w_62_37# s0 0.13fF
C603 enable_0/en a1 0.35fF
C604 4bitadder_1/XOR_1/out 4bitadder_1/XOR_1/w_62_37# 0.02fF
C605 enable_2/en enable_2/a0 0.17fF
C606 a1out_1 a2out_1 7.75fF
C607 comparator_0/t7 comparator_0/t6 0.27fF
C608 comparator_0/4input_AND_1/not_0/in comparator_0/a2xnorb2 0.18fF
C609 comparator_0/xnor_3/XOR_0/w_62_37# comparator_0/xnor_3/not_0/in 0.02fF
C610 b3out_0 4bitadder_0/XOR_3/w_n34_n1# 0.11fF
C611 4bitadder_0/fulladder_2/XOR_0/w_16_n1# vdd 0.02fF
C612 4bitadder_1/fulladder_2/XOR_1/w_62_n20# 4bitadder_1/fulladder_2/XOR_1/abar 0.02fF
C613 4bitadder_0/XOR_3/out gnd 0.42fF
C614 4bitadder_0/fulladder_1/and_0/w_n43_8# 4bitadder_0/fulladder_1/axorb 0.09fF
C615 4bitadder_0/fulladder_2/XOR_0/w_62_n20# 4bitadder_0/fulladder_2/XOR_0/abar 0.02fF
C616 enable_1/en a0 0.24fF
C617 4bitadder_1/fulladder_0/axorb gnd 0.09fF
C618 comparator_0/xnor_0/XOR_0/w_16_n1# comparator_0/b3 0.11fF
C619 4bitadder_0/b0xorM 4bitadder_0/XOR_0/w_62_37# 0.02fF
C620 enable_0/en enable_0/and_3/w_n43_8# 0.09fF
C621 enable_0/and_1/w_26_9# enable_0/and_1/a_n26_14# 0.09fF
C622 vdd 4bitadder_1/fulladder_2/and_0/w_n43_8# 0.07fF
C623 4bitadder_1/c1 4bitadder_1/fulladder_1/XOR_1/w_62_37# 0.13fF
C624 comparator_0/b1bar vdd 0.20fF
C625 enable_2/and_5/a_n26_14# enable_2/and_5/w_26_9# 0.09fF
C626 4bitadder_0/XOR_2/w_62_37# s0 0.13fF
C627 enable_1/and_7/a_n26_14# b3 0.31fF
C628 comparator_0/b3 comparator_0/xnor_0/XOR_0/abar 0.30fF
C629 4bitadder_0/c3 4bitadder_0/fulladder_3/XOR_1/w_62_37# 0.13fF
C630 a2 enable_3/and_2/a_n26_14# 0.31fF
C631 4bitadder_1/c1 s1_sub 0.04fF
C632 vdd comparator_0/xnor_0/XOR_0/w_n34_n1# 0.02fF
C633 4bitadder_1/fulladder_3/XOR_0/w_62_37# 4bitadder_1/XOR_3/out 0.13fF
C634 enable_0/and_1/w_n43_8# vdd 0.07fF
C635 enable_3/and_1/w_n43_8# enable_3/and_1/a_n26_14# 0.02fF
C636 b1out_1 4bitadder_1/XOR_1/abar 0.13fF
C637 a2out_3 vdd 0.12fF
C638 comparator_0/a1bar comparator_0/not_5/w_n2_10# 0.03fF
C639 vdd 4bitadder_1/fulladder_3/or_0/a 0.14fF
C640 4bitadder_1/fulladder_0/XOR_1/bbar s0 0.02fF
C641 4bitadder_1/fulladder_0/axorb 4bitadder_1/fulladder_0/XOR_1/abar 0.13fF
C642 4bitadder_1/fulladder_0/and_0/a_n26_14# s0 0.10fF
C643 a2out_2 comparator_0/3input_AND_0/w_32_n21# 0.16fF
C644 comparator_0/b3 gnd 0.83fF
C645 4bitadder_0/c3 s3_add 0.04fF
C646 enable_1/and_3/w_n43_8# enable_1/and_3/a_n26_14# 0.02fF
C647 4bitadder_1/fulladder_2/and_0/a_n26_14# 4bitadder_1/fulladder_2/and_0/w_n43_8# 0.02fF
C648 comparator_0/b3 comparator_0/not_3/w_n2_10# 0.09fF
C649 4bitadder_0/fulladder_3/XOR_0/w_62_37# 4bitadder_0/XOR_3/out 0.13fF
C650 4bitadder_1/fulladder_0/XOR_0/abar 4bitadder_1/fulladder_0/XOR_0/w_n34_n1# 0.03fF
C651 enable_3/and_5/w_26_9# b1out_3 0.03fF
C652 4bitadder_1/fulladder_0/XOR_0/w_62_n20# 4bitadder_1/fulladder_0/XOR_0/abar 0.02fF
C653 enable_2/and_4/w_26_9# vdd 0.03fF
C654 enable_2/and_0/w_n43_8# vdd 0.07fF
C655 comparator_0/4input_OR_0/w_n58_n43# comparator_0/t7 0.13fF
C656 4bitadder_1/XOR_1/w_62_37# s0 0.13fF
C657 4bitadder_0/XOR_0/w_16_n1# s0 0.11fF
C658 enable_0/and_4/w_26_9# vdd 0.03fF
C659 vdd comparator_0/5input_AND_0/w_31_n55# 0.06fF
C660 b1 a1 0.28fF
C661 enable_0/and_0/a_n26_14# a0 0.31fF
C662 vdd enable_0/and_5/w_n43_8# 0.07fF
C663 b0out_0 gnd 0.15fF
C664 4bitadder_1/fulladder_0/axorb 4bitadder_1/fulladder_0/XOR_0/w_62_37# 0.02fF
C665 b1out_0 4bitadder_0/XOR_1/w_n34_n1# 0.11fF
C666 4bitadder_0/fulladder_1/and_1/w_n43_8# vdd 0.07fF
C667 gnd 4bitadder_1/fulladder_2/XOR_0/abar 0.15fF
C668 4bitadder_0/fulladder_0/XOR_0/abar a0out_0 0.13fF
C669 enable_0/en decoder_0/and_0/w_26_9# 0.03fF
C670 a2out_2 boout_2 0.51fF
C671 b2out_2 a0out_2 0.42fF
C672 gnd b2out_1 0.92fF
C673 enable_3/and_0/w_n43_8# enable_3/en 0.09fF
C674 4bitadder_1/XOR_2/out s0 0.19fF
C675 comparator_0/b3 comparator_0/and_1/w_n43_8# 0.09fF
C676 a1out_2 gnd 0.83fF
C677 4bitadder_1/XOR_2/w_62_37# b2out_1 0.02fF
C678 4bitadder_1/fulladder_3/axorb 4bitadder_1/fulladder_3/XOR_0/w_62_n20# 0.04fF
C679 vdd comparator_0/a3bar 0.04fF
C680 comparator_0/4input_OR_1/y gnd 0.03fF
C681 vdd 4bitadder_1/XOR_1/w_n34_n1# 0.02fF
C682 vdd b1out_2 1.29fF
C683 comparator_0/3input_AND_1/w_69_n71# comparator_0/a3xnorb3 0.16fF
C684 a3out_1 b3out_1 0.20fF
C685 vdd 4bitadder_1/fulladder_1/or_0/a 0.14fF
C686 a3out_2 comparator_0/b3bar 3.31fF
C687 a1out_2 comparator_0/4input_AND_1/w_n47_52# 0.16fF
C688 enable_3/and_1/w_26_9# vdd 0.03fF
C689 a0 b0 0.37fF
C690 vdd 4bitadder_1/c1 0.12fF
C691 comparator_0/xnor_2/XOR_0/w_62_37# a1out_2 0.02fF
C692 enable_0/and_7/w_n43_8# vdd 0.07fF
C693 4bitadder_0/fulladder_1/and_1/w_26_9# 4bitadder_0/fulladder_1/and_1/a_n26_14# 0.09fF
C694 4bitadder_0/fulladder_1/XOR_0/w_n34_n1# vdd 0.02fF
C695 4bitadder_1/XOR_2/w_62_n20# 4bitadder_1/XOR_2/bbar 0.13fF
C696 4bitadder_1/fulladder_2/and_0/w_26_9# 4bitadder_1/fulladder_2/or_0/a 0.03fF
C697 vdd comparator_0/and_1/w_26_9# 0.03fF
C698 a1out_1 gnd 0.92fF
C699 comparator_0/4input_OR_1/w_n58_n43# comparator_0/t4 0.13fF
C700 4bitadder_0/fulladder_0/XOR_1/w_62_n20# 4bitadder_0/fulladder_0/XOR_1/abar 0.02fF
C701 enable_3/and_0/w_26_9# vdd 0.03fF
C702 vdd decoder_0/and_3/w_n43_8# 0.07fF
C703 comparator_0/t4 comparator_0/5input_AND_1/not_0/w_n2_10# 0.03fF
C704 comparator_0/xnor_2/XOR_0/w_62_n20# comparator_0/xnor_2/XOR_0/bbar 0.13fF
C705 4bitadder_0/XOR_2/w_62_n20# 4bitadder_0/XOR_2/bbar 0.13fF
C706 enable_3/and_1/w_26_9# a1out_3 0.03fF
C707 b1out_3 gnd 0.25fF
C708 enable_1/and_6/w_26_9# b2out_1 0.03fF
C709 4bitadder_1/fulladder_0/and_1/a_n26_14# 4bitadder_1/fulladder_0/and_1/w_26_9# 0.09fF
C710 vdd comparator_0/4input_AND_2/w_n47_52# 0.02fF
C711 comparator_0/4input_OR_1/y comparator_0/4input_OR_1/w_n58_n43# 0.02fF
C712 enable_1/and_0/a_n26_14# enable_1/and_0/w_26_9# 0.09fF
C713 4bitadder_1/b0xorM s0 0.26fF
C714 comparator_0/a0xnorb0 gnd 0.36fF
C715 4bitadder_1/fulladder_0/XOR_1/bbar 4bitadder_1/fulladder_0/XOR_1/w_62_n20# 0.13fF
C716 comparator_0/t5 gnd 0.34fF
C717 a0 enable_2/a0 0.05fF
C718 4bitadder_1/XOR_1/w_62_37# b1out_1 0.02fF
C719 comparator_0/4input_AND_2/not_0/in comparator_0/a3xnorb3 0.18fF
C720 a1 a2 0.40fF
C721 enable_2/and_2/w_26_9# enable_2/and_2/a_n26_14# 0.09fF
C722 enable_0/en a3 0.37fF
C723 vdd 4bitadder_1/fulladder_0/or_0/w_n48_101# 0.05fF
C724 4bitadder_0/c1 a1out_0 0.35fF
C725 b1out_0 a2out_0 0.14fF
C726 4bitadder_1/fulladder_0/or_0/a_n15_32# 4bitadder_1/fulladder_0/or_0/b 0.19fF
C727 comparator_0/a1bar comparator_0/a3xnorb3 0.36fF
C728 4bitadder_0/c3 4bitadder_0/fulladder_2/or_0/w_58_101# 0.02fF
C729 comparator_0/4input_OR_1/w_n58_n43# comparator_0/t3 0.13fF
C730 decoder_0/and_0/w_n43_8# decoder_0/and_2/a 0.09fF
C731 comparator_0/3input_AND_0/not_0/in comparator_0/a3xnorb3 0.19fF
C732 4bitadder_0/XOR_1/bbar s0 0.02fF
C733 enable_0/and_2/w_26_9# enable_0/and_2/a_n26_14# 0.09fF
C734 4bitadder_0/fulladder_2/and_0/w_n43_8# 4bitadder_0/c2 0.09fF
C735 a1 vdd 0.42fF
C736 vdd 4bitadder_1/fulladder_1/or_0/w_n48_101# 0.05fF
C737 vdd comparator_0/3input_AND_0/not_0/w_n2_10# 0.18fF
C738 4bitadder_1/fulladder_3/XOR_0/w_62_n20# 4bitadder_1/fulladder_3/XOR_0/bbar 0.13fF
C739 comparator_0/4input_AND_2/not_0/w_n2_10# comparator_0/4input_AND_2/not_0/in 0.09fF
C740 out0 AND_Block_0/and_0/w_26_9# 0.03fF
C741 b1out_0 enable_0/and_5/w_26_9# 0.03fF
C742 4bitadder_1/c1 4bitadder_1/XOR_1/out 0.37fF
C743 a1out_2 comparator_0/a2xnorb2 0.61fF
C744 4bitadder_0/fulladder_2/axorb 4bitadder_0/fulladder_2/XOR_1/w_62_37# 0.02fF
C745 4bitadder_0/fulladder_1/or_0/w_n48_101# vdd 0.05fF
C746 enable_2/and_3/w_n43_8# vdd 0.07fF
C747 comparator_0/xnor_0/not_0/w_n2_10# comparator_0/xnor_0/not_0/in 0.09fF
C748 4bitadder_0/fulladder_3/XOR_0/w_62_n20# 4bitadder_0/fulladder_3/XOR_0/bbar 0.13fF
C749 a3 enable_3/and_3/a_n26_14# 0.31fF
C750 b1out_0 a3out_0 0.12fF
C751 enable_0/and_3/w_n43_8# vdd 0.07fF
C752 4bitadder_0/XOR_3/abar gnd 0.20fF
C753 4bitadder_0/fulladder_0/or_0/a 4bitadder_0/fulladder_0/or_0/w_n48_101# 0.12fF
C754 b2 gnd 0.30fF
C755 comparator_0/4input_AND_2/not_0/in comparator_0/4input_AND_2/w_29_n46# 0.02fF
C756 decoder_0/and_3/w_26_9# decoder_0/and_3/a_n26_14# 0.09fF
C757 vdd a3out_1 0.15fF
C758 enable_1/and_4/w_n43_8# enable_1/and_4/a_n26_14# 0.02fF
C759 enable_1/en a1 0.28fF
C760 vdd a2out_2 1.48fF
C761 comparator_0/xnor_0/not_0/w_n2_10# vdd 0.18fF
C762 4bitadder_0/fulladder_1/or_0/w_n48_101# 4bitadder_0/fulladder_1/or_0/b 0.12fF
C763 enable_3/en enable_3/and_3/w_n43_8# 0.09fF
C764 enable_1/and_6/w_n43_8# b2 0.09fF
C765 4bitadder_1/XOR_0/bbar s0 0.02fF
C766 4bitadder_1/fulladder_1/or_0/w_n48_101# 4bitadder_1/fulladder_1/or_0/b 0.12fF
C767 comparator_0/a0xnorb0 comparator_0/a2xnorb2 0.36fF
C768 comparator_0/xnor_1/XOR_0/abar gnd 0.14fF
C769 enable_3/and_6/a_n26_14# enable_3/and_6/w_n43_8# 0.02fF
C770 a3out_3 b3out_3 0.29fF
C771 enable_3/and_6/w_26_9# b2out_3 0.03fF
C772 a3out_1 b0out_1 0.13fF
C773 4bitadder_1/fulladder_2/and_1/w_n43_8# 4bitadder_1/XOR_2/out 0.09fF
C774 4bitadder_0/c3 gnd 0.91fF
C775 b1 a3 0.28fF
C776 vdd 4bitadder_1/fulladder_2/XOR_1/w_16_n1# 0.02fF
C777 enable_2/and_0/w_n43_8# enable_2/a0 0.09fF
C778 enable_2/b1 gnd 0.07fF
C779 comparator_0/xnor_3/XOR_0/w_62_n20# comparator_0/xnor_3/XOR_0/bbar 0.13fF
C780 enable_3/and_6/a_n26_14# enable_3/and_6/w_26_9# 0.09fF
C781 4bitadder_1/XOR_1/w_16_n1# 4bitadder_1/XOR_1/bbar 0.03fF
C782 4bitadder_1/b0xorM 4bitadder_1/XOR_0/w_62_n20# 0.04fF
C783 comparator_0/t6 comparator_0/3input_AND_0/not_0/w_n2_10# 0.03fF
C784 4bitadder_0/fulladder_0/axorb 4bitadder_0/fulladder_0/XOR_0/w_62_37# 0.02fF
C785 vdd comparator_0/not_7/w_n2_10# 0.26fF
C786 b1out_0 vdd 0.13fF
C787 4bitadder_1/fulladder_3/axorb 4bitadder_1/fulladder_3/XOR_1/w_n34_n1# 0.11fF
C788 comparator_0/4input_OR_1/NOT_0/w_n2_10# comparator_0/4input_OR_1/y 0.09fF
C789 4bitadder_0/XOR_1/w_16_n1# 4bitadder_0/XOR_1/bbar 0.03fF
C790 enable_0/and_5/a_n26_14# enable_0/and_5/w_n43_8# 0.02fF
C791 4bitadder_1/fulladder_1/axorb 4bitadder_1/fulladder_1/XOR_1/w_62_37# 0.02fF
C792 comparator_0/5input_AND_1/not_0/in comparator_0/5input_AND_1/w_31_n55# 0.03fF
C793 enable_2/and_5/w_26_9# vdd 0.03fF
C794 vdd decoder_0/and_0/w_26_9# 0.03fF
C795 vdd 4bitadder_1/fulladder_3/or_0/w_58_101# 0.05fF
C796 4bitadder_0/b0xorM 4bitadder_0/XOR_0/w_62_n20# 0.04fF
C797 AND_Block_0/and_1/w_n43_8# AND_Block_0/and_1/a_n26_14# 0.02fF
C798 s0 decoder_0/and_3/w_n43_8# 0.09fF
C799 4bitadder_0/fulladder_2/XOR_1/abar gnd 0.15fF
C800 enable_0/and_6/w_n43_8# enable_0/and_6/a_n26_14# 0.02fF
C801 4bitadder_0/XOR_2/out a2out_0 1.88fF
C802 4bitadder_0/fulladder_2/and_1/w_26_9# 4bitadder_0/fulladder_2/or_0/b 0.03fF
C803 4bitadder_1/fulladder_2/axorb 4bitadder_1/XOR_2/out 0.13fF
C804 4bitadder_1/fulladder_1/or_0/w_n48_101# 4bitadder_1/fulladder_1/or_0/a_n15_32# 0.05fF
C805 4bitadder_0/fulladder_3/XOR_1/abar gnd 0.15fF
C806 enable_2/and_3/w_26_9# enable_2/and_3/a_n26_14# 0.09fF
C807 a2 a3 0.21fF
C808 a1 b0 0.37fF
C809 vdd comparator_0/3input_AND_0/w_n14_24# 0.03fF
C810 enable_2/a2 gnd 0.07fF
C811 4bitadder_1/XOR_1/w_n34_n1# b1out_1 0.11fF
C812 comparator_0/4input_OR_0/NOT_0/w_n2_10# comparator_0/4input_OR_0/y 0.09fF
C813 4bitadder_1/XOR_0/bbar 4bitadder_1/XOR_0/w_62_n20# 0.13fF
C814 comparator_0/3input_AND_1/not_0/in comparator_0/3input_AND_1/w_32_n21# 0.02fF
C815 enable_0/and_3/w_26_9# enable_0/and_3/a_n26_14# 0.09fF
C816 a3 vdd 0.44fF
C817 4bitadder_1/XOR_3/out a3out_1 2.13fF
C818 4bitadder_1/fulladder_3/and_1/w_26_9# 4bitadder_1/fulladder_3/or_0/b 0.03fF
C819 comparator_0/b3 boout_2 0.36fF
C820 4bitadder_0/fulladder_3/or_0/w_n48_101# 4bitadder_0/fulladder_3/or_0/b 0.12fF
C821 4bitadder_1/c1 4bitadder_1/fulladder_1/and_0/w_n43_8# 0.09fF
C822 enable_3/and_1/w_n43_8# vdd 0.07fF
C823 4bitadder_1/fulladder_0/XOR_0/w_62_n20# 4bitadder_1/fulladder_0/axorb 0.04fF
C824 comparator_0/b2bar comparator_0/a3xnorb3 0.38fF
C825 comparator_0/xnor_1/XOR_0/w_62_37# comparator_0/xnor_1/not_0/in 0.02fF
C826 b0 enable_3/and_4/a_n26_14# 0.31fF
C827 4bitadder_0/XOR_3/out a3out_0 2.19fF
C828 4bitadder_0/fulladder_3/and_1/w_26_9# 4bitadder_0/fulladder_3/or_0/b 0.03fF
C829 4bitadder_0/fulladder_0/and_1/w_n43_8# 4bitadder_0/b0xorM 0.09fF
C830 4bitadder_1/fulladder_2/XOR_0/w_62_37# a2out_1 0.02fF
C831 4bitadder_0/fulladder_1/and_0/w_n43_8# vdd 0.07fF
C832 vdd 4bitadder_1/fulladder_2/and_1/w_26_9# 0.03fF
C833 vdd 4bitadder_1/fulladder_1/axorb 0.15fF
C834 enable_3/and_6/w_n43_8# vdd 0.07fF
C835 4bitadder_1/fulladder_2/axorb 4bitadder_1/fulladder_2/and_0/w_n43_8# 0.09fF
C836 b2out_2 comparator_0/xnor_1/XOR_0/bbar 0.02fF
C837 comparator_0/4input_OR_1/w_n58_n43# comparator_0/t2 0.13fF
C838 4bitadder_0/XOR_0/bbar 4bitadder_0/XOR_0/w_62_n20# 0.13fF
C839 enable_2/and_1/w_n43_8# enable_2/en 0.09fF
C840 enable_2/and_7/w_26_9# b3out_2 0.03fF
C841 enable_1/en a3 0.28fF
C842 gnd 4bitadder_1/fulladder_2/or_0/b 0.37fF
C843 enable_3/en gnd 0.13fF
C844 4bitadder_1/fulladder_2/XOR_0/bbar 4bitadder_1/XOR_2/out 0.02fF
C845 4bitadder_1/fulladder_0/or_0/b gnd 0.37fF
C846 4bitadder_0/fulladder_0/or_0/w_n48_101# 4bitadder_0/fulladder_0/or_0/b 0.12fF
C847 4bitadder_1/XOR_2/out 4bitadder_1/XOR_2/w_62_n20# 0.04fF
C848 4bitadder_0/fulladder_0/or_0/w_n48_101# 4bitadder_0/fulladder_0/or_0/a_n15_32# 0.05fF
C849 vdd comparator_0/not_6/w_n2_10# 0.18fF
C850 enable_3/and_6/w_26_9# vdd 0.03fF
C851 4bitadder_0/fulladder_0/and_0/a_n26_14# s0 0.10fF
C852 enable_2/and_6/w_26_9# b2out_2 0.03fF
C853 b2out_3 b1out_3 29.73fF
C854 AND_Block_0/and_1/w_26_9# AND_Block_0/and_1/a_n26_14# 0.09fF
C855 enable_2/and_6/w_n43_8# enable_2/en 0.09fF
C856 enable_2/and_5/w_n43_8# enable_2/and_5/a_n26_14# 0.02fF
C857 a1out_2 boout_2 0.64fF
C858 b1out_2 a0out_2 1.11fF
C859 b0out_0 a2out_0 0.12fF
C860 comparator_0/3input_AND_0/not_0/in comparator_0/3input_AND_0/w_69_n71# 0.02fF
C861 comparator_0/not_6/w_n2_10# comparator_0/a2bar 0.03fF
C862 4bitadder_0/fulladder_0/and_0/w_26_9# 4bitadder_0/fulladder_0/and_0/a_n26_14# 0.09fF
C863 b1out_0 s0 13.84fF
C864 enable_2/and_5/a_n26_14# enable_2/b1 0.31fF
C865 4bitadder_1/XOR_1/out 4bitadder_1/fulladder_1/XOR_0/bbar 0.02fF
C866 b2out_0 4bitadder_0/XOR_2/w_n34_n1# 0.11fF
C867 4bitadder_1/fulladder_2/XOR_1/w_n34_n1# 4bitadder_1/fulladder_2/XOR_1/abar 0.03fF
C868 4bitadder_1/fulladder_2/XOR_1/w_16_n1# 4bitadder_1/fulladder_2/XOR_1/bbar 0.03fF
C869 4bitadder_1/fulladder_2/XOR_1/w_62_n20# s2_sub 0.04fF
C870 comparator_0/xnor_0/XOR_0/w_62_37# comparator_0/b3 0.13fF
C871 enable_1/and_5/a_n26_14# b1 0.31fF
C872 4bitadder_1/fulladder_0/axorb vdd 0.15fF
C873 4bitadder_0/fulladder_2/axorb gnd 0.09fF
C874 4bitadder_0/XOR_0/w_62_37# s0 0.13fF
C875 a1out_1 b3out_1 0.24fF
C876 b0out_0 a3out_0 0.12fF
C877 4bitadder_0/fulladder_2/and_0/w_26_9# 4bitadder_0/fulladder_2/and_0/a_n26_14# 0.09fF
C878 enable_0/en b2 0.38fF
C879 a3out_1 b1out_1 0.18fF
C880 enable_3/en decoder_0/and_3/w_26_9# 0.03fF
C881 4bitadder_1/fulladder_1/axorb 4bitadder_1/XOR_1/out 0.13fF
C882 comparator_0/b3 comparator_0/xnor_0/not_0/in 0.13fF
C883 a3out_2 comparator_0/xnor_0/XOR_0/abar 0.13fF
C884 4bitadder_0/fulladder_2/XOR_1/w_62_37# s2_add 0.02fF
C885 a3out_2 gnd 0.76fF
C886 vdd comparator_0/b3 0.82fF
C887 enable_1/and_3/w_26_9# vdd 0.03fF
C888 a3 b0 0.37fF
C889 4bitadder_1/fulladder_2/or_0/a_n15_32# 4bitadder_1/fulladder_2/or_0/w_n48_101# 0.05fF
C890 enable_2/and_4/w_26_9# enable_2/and_4/a_n26_14# 0.09fF
C891 b2 enable_3/and_6/a_n26_14# 0.31fF
C892 comparator_0/5input_AND_0/not_0/in comparator_0/5input_AND_0/w_106_n113# 0.03fF
C893 vdd 4bitadder_1/fulladder_2/XOR_0/w_16_n1# 0.02fF
C894 vdd comparator_0/5input_AND_0/w_n37_15# 0.05fF
C895 enable_1/and_0/w_n43_8# a0 0.09fF
C896 enable_0/and_4/w_26_9# enable_0/and_4/a_n26_14# 0.09fF
C897 4bitadder_1/XOR_1/w_62_n20# 4bitadder_1/XOR_1/bbar 0.13fF
C898 comparator_0/5input_AND_1/not_0/in gnd 0.10fF
C899 comparator_0/5input_AND_0/not_0/in comparator_0/a3xnorb3 0.23fF
C900 b0out_0 vdd 0.13fF
C901 4bitadder_0/fulladder_0/XOR_0/bbar 4bitadder_0/b0xorM 0.02fF
C902 4bitadder_0/fulladder_0/axorb 4bitadder_0/fulladder_0/XOR_0/w_62_n20# 0.04fF
C903 4bitadder_1/fulladder_3/XOR_1/w_62_37# s3_sub 0.02fF
C904 4bitadder_0/fulladder_0/XOR_1/w_n34_n1# vdd 0.02fF
C905 4bitadder_1/fulladder_2/XOR_0/w_62_n20# 4bitadder_1/fulladder_2/XOR_0/abar 0.02fF
C906 a2out_2 a0out_2 0.55fF
C907 vdd comparator_0/t4 0.04fF
C908 a0out_3 gnd 0.11fF
C909 vdd b2out_1 0.05fF
C910 4bitadder_0/XOR_1/out gnd 0.42fF
C911 vdd 4bitadder_1/XOR_1/w_16_n1# 0.02fF
C912 vdd a1out_2 1.25fF
C913 4bitadder_0/XOR_1/w_62_n20# 4bitadder_0/XOR_1/bbar 0.13fF
C914 4bitadder_0/fulladder_3/XOR_1/w_62_37# s3_add 0.02fF
C915 b2 b1 0.23fF
C916 4bitadder_1/XOR_3/out 4bitadder_1/XOR_3/w_62_n20# 0.04fF
C917 comparator_0/a1xnorb1 comparator_0/5input_AND_0/not_0/in 0.23fF
C918 out3 AND_Block_0/and_3/w_26_9# 0.03fF
C919 gnd 4bitadder_1/XOR_2/abar 0.13fF
C920 4bitadder_0/fulladder_2/XOR_0/abar gnd 0.15fF
C921 b3out_3 gnd 0.24fF
C922 gnd 4bitadder_1/XOR_0/abar 0.15fF
C923 comparator_0/xnor_2/XOR_0/abar gnd 0.14fF
C924 4bitadder_0/XOR_3/out 4bitadder_0/XOR_3/w_62_n20# 0.04fF
C925 4bitadder_0/fulladder_1/and_1/w_n43_8# a1out_0 0.09fF
C926 4bitadder_0/fulladder_0/XOR_0/w_n34_n1# vdd 0.02fF
C927 vdd comparator_0/xnor_3/XOR_0/w_n34_n1# 0.02fF
C928 4bitadder_0/XOR_2/out s0 0.19fF
C929 AND_Block_0/and_0/w_n43_8# b0out_3 0.09fF
C930 vdd a1out_1 0.33fF
C931 comparator_0/a1xnorb1 comparator_0/5input_AND_0/w_106_n113# 0.17fF
C932 4bitadder_0/fulladder_0/XOR_1/w_n34_n1# 4bitadder_0/fulladder_0/XOR_1/abar 0.03fF
C933 4bitadder_0/fulladder_0/XOR_1/w_16_n1# 4bitadder_0/fulladder_0/XOR_1/bbar 0.03fF
C934 4bitadder_0/fulladder_0/XOR_1/w_62_n20# s0_add 0.04fF
C935 comparator_0/5input_AND_1/not_0/in comparator_0/5input_AND_1/not_0/w_n2_10# 0.09fF
C936 4bitadder_0/fulladder_1/XOR_0/w_16_n1# vdd 0.02fF
C937 a3out_2 comparator_0/a2xnorb2 0.15fF
C938 b1out_3 vdd 0.12fF
C939 vdd comparator_0/t3 0.04fF
C940 comparator_0/4input_AND_0/not_0/w_n2_10# equal 0.03fF
C941 comparator_0/a1xnorb1 comparator_0/a3xnorb3 1.11fF
C942 comparator_0/b3bar gnd 0.27fF
C943 comparator_0/not_3/w_n2_10# comparator_0/b3bar 0.03fF
C944 b2out_0 4bitadder_0/XOR_1/abar 1.51fF
C945 vdd comparator_0/a0xnorb0 0.04fF
C946 4bitadder_0/fulladder_3/XOR_0/abar gnd 0.15fF
C947 4bitadder_0/fulladder_1/XOR_0/w_n34_n1# a1out_0 0.11fF
C948 b1 enable_2/b1 0.08fF
C949 a1out_1 b0out_1 0.11fF
C950 comparator_0/a0bar comparator_0/a2xnorb2 0.41fF
C951 comparator_0/4input_AND_0/not_0/in comparator_0/4input_AND_0/w_68_n95# 0.02fF
C952 enable_2/and_2/w_n43_8# enable_2/a2 0.09fF
C953 4bitadder_0/XOR_3/out s0 0.16fF
C954 4bitadder_0/fulladder_1/axorb 4bitadder_0/XOR_1/out 0.13fF
C955 4bitadder_0/fulladder_1/XOR_0/w_62_37# a1out_0 0.02fF
C956 4bitadder_1/fulladder_0/axorb s0 0.54fF
C957 a1out_3 b1out_3 2.06fF
C958 enable_2/and_3/w_26_9# a3out_2 0.03fF
C959 b1out_2 comparator_0/4input_AND_2/not_0/in 0.18fF
C960 4bitadder_0/XOR_1/out 4bitadder_0/XOR_1/w_62_37# 0.02fF
C961 enable_1/and_2/w_n43_8# a2 0.09fF
C962 b3 enable_2/en 0.22fF
C963 comparator_0/a1bar b1out_2 0.44fF
C964 comparator_0/5input_AND_1/not_0/in comparator_0/a2xnorb2 0.23fF
C965 comparator_0/xnor_2/not_0/w_n2_10# comparator_0/xnor_2/not_0/in 0.09fF
C966 4bitadder_0/c3 a3out_0 0.36fF
C967 enable_0/and_6/w_26_9# vdd 0.03fF
C968 b2 a2 0.21fF
C969 4bitadder_0/XOR_3/w_16_n1# vdd 0.02fF
C970 enable_1/and_2/w_n43_8# vdd 0.07fF
C971 4bitadder_1/fulladder_1/axorb 4bitadder_1/fulladder_1/and_0/w_n43_8# 0.09fF
C972 b2out_0 gnd 1.03fF
C973 4bitadder_1/fulladder_2/axorb 4bitadder_1/fulladder_2/XOR_1/abar 0.13fF
C974 a1out_1 4bitadder_1/XOR_1/out 1.87fF
C975 4bitadder_1/b0xorM a0_out1 1.79fF
C976 comparator_0/4input_AND_2/not_0/in comparator_0/4input_AND_2/w_n47_52# 0.02fF
C977 a3out_3 gnd 0.14fF
C978 decoder_0/and_3/w_n43_8# s1 0.09fF
C979 enable_0/and_0/w_n43_8# a0 0.09fF
C980 b2 vdd 0.45fF
C981 comparator_0/a1bar comparator_0/4input_AND_2/w_n47_52# 0.16fF
C982 gnd 4bitadder_1/fulladder_2/or_0/a 0.01fF
C983 vdd comparator_0/xnor_1/XOR_0/w_16_n1# 0.02fF
C984 4bitadder_0/fulladder_0/XOR_0/w_62_n20# 4bitadder_0/fulladder_0/XOR_0/abar 0.02fF
C985 comparator_0/4input_OR_0/y gnd 0.03fF
C986 4bitadder_0/fulladder_0/and_1/w_n43_8# vdd 0.07fF
C987 enable_1/en enable_1/and_2/w_n43_8# 0.09fF
C988 enable_1/and_7/w_26_9# b3out_1 0.03fF
C989 4bitadder_1/fulladder_3/or_0/a_n15_32# 4bitadder_1/fulladder_3/or_0/b 0.19fF
C990 comparator_0/b3bar comparator_0/a2xnorb2 0.12fF
C991 comparator_0/t5 comparator_0/t6 0.21fF
C992 comparator_0/xnor_1/not_0/in gnd 0.03fF
C993 b1 enable_2/a2 0.09fF
C994 enable_2/and_5/w_n43_8# vdd 0.07fF
C995 b0out_0 s0 0.15fF
C996 4bitadder_0/c3 vdd 0.12fF
C997 enable_3/and_0/a_n26_14# a0 0.31fF
C998 enable_1/en b2 0.28fF
C999 s0 b2out_1 0.35fF
C1000 b2out_2 comparator_0/a3xnorb3 0.19fF
C1001 4bitadder_0/fulladder_0/axorb 4bitadder_0/fulladder_0/XOR_1/w_n34_n1# 0.11fF
C1002 4bitadder_1/XOR_1/w_16_n1# s0 0.11fF
C1003 comparator_0/a0bar comparator_0/5input_AND_1/w_n37_15# 0.17fF
C1004 vdd comparator_0/not_4/w_n2_10# 0.26fF
C1005 enable_2/b1 vdd 0.12fF
C1006 vdd s2_sub 0.19fF
C1007 comparator_0/3input_AND_0/not_0/in comparator_0/3input_AND_0/not_0/w_n2_10# 0.09fF
C1008 4bitadder_0/fulladder_0/XOR_1/bbar s0 0.02fF
C1009 4bitadder_0/fulladder_2/XOR_1/w_16_n1# vdd 0.02fF
C1010 4bitadder_0/fulladder_1/XOR_0/abar 4bitadder_0/XOR_1/out 0.25fF
C1011 b2out_2 comparator_0/a1xnorb1 0.27fF
C1012 enable_3/and_5/w_n43_8# enable_3/en 0.09fF
C1013 gnd 4bitadder_1/fulladder_3/axorb 0.09fF
C1014 vdd 4bitadder_1/fulladder_1/and_1/w_26_9# 0.03fF
C1015 enable_2/en decoder_0/and_2/w_26_9# 0.03fF
C1016 a1out_1 s0 0.21fF
C1017 comparator_0/5input_AND_1/not_0/in comparator_0/5input_AND_1/w_n37_15# 0.05fF
C1018 vdd comparator_0/5input_AND_1/w_106_n113# 0.04fF
C1019 4bitadder_0/fulladder_1/and_0/w_26_9# 4bitadder_0/fulladder_1/and_0/a_n26_14# 0.09fF
C1020 4bitadder_1/XOR_3/w_n34_n1# b3out_1 0.11fF
C1021 4bitadder_1/c3 4bitadder_1/fulladder_3/XOR_1/bbar 0.02fF
C1022 enable_3/en b1 0.25fF
C1023 4bitadder_0/fulladder_2/and_1/w_n43_8# 4bitadder_0/fulladder_2/and_1/a_n26_14# 0.02fF
C1024 a2out_2 comparator_0/3input_AND_0/not_0/in 0.19fF
C1025 comparator_0/4input_OR_0/w_n58_n43# comparator_0/t5 0.13fF
C1026 4bitadder_0/fulladder_3/XOR_1/w_16_n1# vdd 0.02fF
C1027 4bitadder_0/fulladder_1/XOR_1/w_62_n20# 4bitadder_0/fulladder_1/XOR_1/bbar 0.13fF
C1028 4bitadder_0/fulladder_0/XOR_0/w_16_n1# 4bitadder_0/fulladder_0/XOR_0/bbar 0.03fF
C1029 4bitadder_1/c2 4bitadder_1/XOR_2/out 0.55fF
C1030 4bitadder_1/XOR_3/w_62_n20# 4bitadder_1/XOR_3/abar 0.02fF
C1031 4bitadder_0/fulladder_3/or_0/w_58_101# vdd 0.05fF
C1032 a2 enable_2/a2 0.11fF
C1033 4bitadder_1/fulladder_0/and_1/a_n26_14# a0_out1 0.10fF
C1034 vdd comparator_0/4input_AND_0/not_0/w_n2_10# 0.18fF
C1035 4bitadder_1/fulladder_1/and_1/w_26_9# 4bitadder_1/fulladder_1/or_0/b 0.03fF
C1036 4bitadder_0/XOR_3/w_62_n20# 4bitadder_0/XOR_3/abar 0.02fF
C1037 AND_Block_0/and_3/a_n26_14# AND_Block_0/and_3/w_n43_8# 0.02fF
C1038 a1 enable_2/and_1/w_n43_8# 0.09fF
C1039 enable_0/and_0/w_26_9# a0out_0 0.03fF
C1040 a0 b3 0.32fF
C1041 enable_1/and_7/w_26_9# vdd 0.03fF
C1042 enable_1/and_3/w_n43_8# a3 0.09fF
C1043 b1out_1 b2out_1 0.26fF
C1044 enable_2/a2 vdd 0.10fF
C1045 4bitadder_1/fulladder_1/XOR_1/w_62_n20# 4bitadder_1/fulladder_1/XOR_1/bbar 0.13fF
C1046 4bitadder_1/fulladder_0/and_1/w_n43_8# vdd 0.07fF
C1047 4bitadder_1/fulladder_0/or_0/a_n15_32# 4bitadder_1/fulladder_0/or_0/w_58_101# 0.13fF
C1048 vdd comparator_0/4input_AND_0/w_29_n46# 0.02fF
C1049 4bitadder_0/c2 4bitadder_0/XOR_2/out 0.55fF
C1050 comparator_0/3input_AND_1/not_0/in gnd 0.21fF
C1051 4bitadder_0/XOR_3/w_16_n1# s0 0.11fF
C1052 4bitadder_0/XOR_0/w_n34_n1# vdd 0.02fF
C1053 out3 gnd 0.01fF
C1054 4bitadder_0/fulladder_2/and_0/a_n26_14# 4bitadder_0/c2 0.10fF
C1055 4bitadder_1/fulladder_0/XOR_0/abar a0_out1 0.13fF
C1056 vdd comparator_0/t2 0.04fF
C1057 4bitadder_1/fulladder_3/and_1/w_n43_8# 4bitadder_1/fulladder_3/and_1/a_n26_14# 0.02fF
C1058 4bitadder_1/fulladder_0/XOR_1/w_16_n1# 4bitadder_1/fulladder_0/XOR_1/bbar 0.03fF
C1059 b2 b0 0.34fF
C1060 a3out_2 boout_2 0.37fF
C1061 comparator_0/b3 a0out_2 0.58fF
C1062 enable_1/and_4/w_n43_8# vdd 0.07fF
C1063 comparator_0/xnor_1/XOR_0/w_n34_n1# a2out_2 0.11fF
C1064 4bitadder_0/XOR_3/abar s0 0.30fF
C1065 decoder_0/and_0/a_n26_14# decoder_0/and_1/b 0.33fF
C1066 comparator_0/3input_AND_0/w_69_n71# comparator_0/a3xnorb3 0.16fF
C1067 4bitadder_0/fulladder_3/and_1/w_n43_8# 4bitadder_0/fulladder_3/and_1/a_n26_14# 0.02fF
C1068 enable_2/and_1/w_26_9# enable_2/and_1/a_n26_14# 0.09fF
C1069 b3out_2 gnd 0.16fF
C1070 comparator_0/4input_AND_1/not_0/in comparator_0/4input_AND_1/w_68_n95# 0.02fF
C1071 comparator_0/a0bar boout_2 0.33fF
C1072 enable_3/en a2 0.25fF
C1073 enable_0/and_7/w_26_9# enable_0/and_7/a_n26_14# 0.09fF
C1074 a0out_2 comparator_0/5input_AND_0/w_n37_15# 0.17fF
C1075 4bitadder_1/c2 4bitadder_1/fulladder_2/and_0/w_n43_8# 0.09fF
C1076 comparator_0/xnor_1/XOR_0/w_62_n20# comparator_0/xnor_1/XOR_0/abar 0.02fF
C1077 gnd a2out_1 1.13fF
C1078 comparator_0/and_1/a_n26_14# gnd 0.02fF
C1079 enable_1/en enable_1/and_4/w_n43_8# 0.09fF
C1080 vdd 4bitadder_1/XOR_3/w_n34_n1# 0.02fF
C1081 boout_2 comparator_0/5input_AND_1/not_0/in 0.23fF
C1082 4bitadder_0/fulladder_2/and_1/w_26_9# vdd 0.03fF
C1083 4bitadder_0/fulladder_2/XOR_0/w_n34_n1# 4bitadder_0/fulladder_2/XOR_0/abar 0.03fF
C1084 enable_3/en vdd 0.68fF
C1085 enable_3/and_0/a_n26_14# enable_3/and_0/w_26_9# 0.09fF
C1086 a1out_2 a0out_2 0.58fF
C1087 comparator_0/5input_AND_0/not_0/in comparator_0/5input_AND_0/not_0/w_n2_10# 0.09fF
C1088 comparator_0/3input_AND_0/not_0/in comparator_0/3input_AND_0/w_n14_24# 0.03fF
C1089 comparator_0/a0xnorb0 comparator_0/4input_AND_0/w_68_n95# 0.16fF
C1090 4bitadder_0/fulladder_2/or_0/b gnd 0.37fF
C1091 4bitadder_0/fulladder_1/XOR_1/abar gnd 0.15fF
C1092 4bitadder_0/fulladder_0/XOR_0/w_n34_n1# 4bitadder_0/fulladder_0/XOR_0/abar 0.03fF
C1093 enable_2/and_7/w_n43_8# vdd 0.07fF
C1094 vdd 4bitadder_1/fulladder_2/and_0/w_26_9# 0.03fF
C1095 4bitadder_0/fulladder_3/or_0/w_n48_101# vdd 0.05fF
C1096 comparator_0/xnor_3/XOR_0/w_n34_n1# a0out_2 0.11fF
C1097 enable_2/and_1/w_26_9# a1out_2 0.03fF
C1098 4bitadder_1/fulladder_0/or_0/b 4bitadder_1/fulladder_0/and_1/w_26_9# 0.03fF
C1099 fc_sub 4bitadder_1/fulladder_3/or_0/w_58_101# 0.02fF
C1100 gnd 4bitadder_1/fulladder_1/XOR_1/abar 0.15fF
C1101 comparator_0/xnor_0/XOR_0/w_62_37# a3out_2 0.02fF
C1102 4bitadder_0/fulladder_3/and_1/w_26_9# vdd 0.03fF
C1103 4bitadder_1/XOR_1/out 4bitadder_1/XOR_1/w_62_n20# 0.04fF
C1104 vdd 4bitadder_1/fulladder_3/or_0/w_n48_101# 0.05fF
C1105 comparator_0/and_1/w_n43_8# comparator_0/and_1/a_n26_14# 0.02fF
C1106 comparator_0/and_1/w_26_9# comparator_0/t1 0.03fF
C1107 4bitadder_0/fulladder_2/axorb vdd 0.15fF
C1108 4bitadder_0/fulladder_3/or_0/b gnd 0.37fF
C1109 4bitadder_0/fulladder_2/XOR_0/abar a2out_0 0.13fF
C1110 enable_1/and_1/a_n26_14# a1 0.31fF
C1111 enable_3/and_7/w_n43_8# enable_3/en 0.09fF
C1112 4bitadder_1/fulladder_2/and_0/a_n26_14# 4bitadder_1/fulladder_2/and_0/w_26_9# 0.09fF
C1113 4bitadder_1/fulladder_0/XOR_0/w_62_n20# 4bitadder_1/fulladder_0/XOR_0/bbar 0.13fF
C1114 comparator_0/xnor_0/XOR_0/w_62_n20# comparator_0/xnor_0/XOR_0/bbar 0.13fF
C1115 4bitadder_0/fulladder_2/or_0/w_n48_101# 4bitadder_0/fulladder_2/or_0/b 0.12fF
C1116 enable_3/and_2/w_n43_8# enable_3/and_2/a_n26_14# 0.02fF
C1117 4bitadder_0/XOR_1/abar gnd 0.23fF
C1118 4bitadder_1/c3 4bitadder_1/fulladder_3/axorb 0.60fF
C1119 comparator_0/b1bar comparator_0/4input_AND_1/w_n8_2# 0.16fF
C1120 4bitadder_0/fulladder_2/XOR_0/w_16_n1# 4bitadder_0/fulladder_2/XOR_0/bbar 0.03fF
C1121 b2out_3 a3out_3 0.13fF
C1122 comparator_0/b1bar comparator_0/a3xnorb3 0.35fF
C1123 vdd a3out_2 0.91fF
C1124 4bitadder_0/fulladder_3/axorb 4bitadder_0/XOR_3/out 0.13fF
C1125 4bitadder_0/c1 4bitadder_0/fulladder_1/XOR_1/bbar 0.02fF
C1126 4bitadder_0/fulladder_1/axorb 4bitadder_0/fulladder_1/XOR_1/abar 0.13fF
C1127 enable_3/and_2/w_26_9# vdd 0.03fF
C1128 enable_1/and_0/w_26_9# vdd 0.03fF
C1129 enable_0/and_7/w_n43_8# b3 0.09fF
C1130 b0 enable_2/a2 0.12fF
C1131 4bitadder_0/fulladder_2/XOR_1/w_62_n20# 4bitadder_0/fulladder_2/XOR_1/abar 0.02fF
C1132 4bitadder_1/fulladder_0/axorb 4bitadder_1/fulladder_0/XOR_1/w_n34_n1# 0.11fF
C1133 decoder_0/and_1/b decoder_0/not_1/w_n2_10# 0.03fF
C1134 a2out_2 comparator_0/b2bar 0.44fF
C1135 comparator_0/xnor_0/XOR_0/abar gnd 0.14fF
C1136 4bitadder_1/fulladder_3/XOR_0/abar a3out_1 0.13fF
C1137 comparator_0/5input_AND_0/not_0/in comparator_0/5input_AND_0/w_31_n55# 0.03fF
C1138 vdd comparator_0/t8 0.04fF
C1139 vdd comparator_0/a0bar 0.30fF
C1140 enable_1/and_4/w_n43_8# b0 0.09fF
C1141 comparator_0/b1bar comparator_0/not_1/w_n2_10# 0.03fF
C1142 vdd 4bitadder_1/fulladder_3/XOR_1/w_n34_n1# 0.02fF
C1143 4bitadder_1/fulladder_1/and_0/a_n26_14# 4bitadder_1/fulladder_1/and_0/w_26_9# 0.09fF
C1144 4bitadder_1/b0xorM 4bitadder_1/fulladder_0/XOR_0/w_16_n1# 0.11fF
C1145 a2out_3 b0out_3 0.16fF
C1146 4bitadder_0/fulladder_3/XOR_0/abar a3out_0 0.13fF
C1147 vdd comparator_0/3input_AND_1/w_32_n21# 0.03fF
C1148 4bitadder_1/fulladder_2/XOR_0/w_n34_n1# 4bitadder_1/fulladder_2/XOR_0/abar 0.03fF
C1149 4bitadder_1/fulladder_2/XOR_0/w_16_n1# 4bitadder_1/fulladder_2/XOR_0/bbar 0.03fF
C1150 b2out_0 a2out_0 0.30fF
C1151 a0out_3 vdd 0.13fF
C1152 vdd 4bitadder_1/XOR_2/w_16_n1# 0.02fF
C1153 vdd comparator_0/4input_AND_1/w_29_n46# 0.02fF
C1154 vdd comparator_0/xnor_2/XOR_0/w_16_n1# 0.02fF
C1155 comparator_0/5input_AND_0/w_31_n55# comparator_0/a3xnorb3 0.21fF
C1156 enable_2/and_7/w_26_9# vdd 0.03fF
C1157 4bitadder_1/fulladder_3/XOR_1/w_62_n20# 4bitadder_1/fulladder_3/XOR_1/abar 0.02fF
C1158 enable_3/en b0 0.25fF
C1159 b3 a1 0.31fF
C1160 comparator_0/xnor_2/not_0/in gnd 0.03fF
C1161 b0out_0 a1out_0 0.11fF
C1162 a0out_3 a1out_3 23.76fF
C1163 gnd 4bitadder_1/fulladder_0/XOR_1/abar 0.15fF
C1164 4bitadder_0/fulladder_3/XOR_1/w_62_n20# 4bitadder_0/fulladder_3/XOR_1/abar 0.02fF
C1165 b2out_0 a3out_0 0.11fF
C1166 comparator_0/xnor_2/XOR_0/w_62_37# comparator_0/xnor_2/not_0/in 0.02fF
C1167 comparator_0/not_4/w_n2_10# a0out_2 0.09fF
C1168 vdd 4bitadder_1/fulladder_0/and_0/w_n43_8# 0.07fF
C1169 b1out_2 comparator_0/a3xnorb3 0.36fF
C1170 4bitadder_0/fulladder_3/XOR_0/w_16_n1# vdd 0.02fF
C1171 a1out_0 4bitadder_0/fulladder_1/and_1/a_n26_14# 0.10fF
C1172 s0 4bitadder_1/XOR_3/bbar 0.02fF
C1173 4bitadder_1/fulladder_1/XOR_0/w_62_n20# 4bitadder_1/fulladder_1/XOR_0/abar 0.02fF
C1174 vdd comparator_0/xnor_3/not_0/w_n2_10# 0.18fF
C1175 4bitadder_1/fulladder_1/XOR_0/w_16_n1# 4bitadder_1/fulladder_1/XOR_0/bbar 0.03fF
C1176 comparator_0/4input_OR_0/NOT_0/w_n2_10# agb 0.03fF
C1177 4bitadder_0/fulladder_1/axorb gnd 0.09fF
C1178 b0out_1 4bitadder_1/XOR_0/abar 0.13fF
C1179 vdd comparator_0/xnor_2/not_0/w_n2_10# 0.18fF
C1180 vdd comparator_0/b3bar 0.04fF
C1181 a0 enable_2/en 0.10fF
C1182 b1out_2 comparator_0/xnor_2/XOR_0/bbar 0.02fF
C1183 comparator_0/a1xnorb1 b1out_2 0.69fF
C1184 comparator_0/t8 comparator_0/t6 0.29fF
C1185 comparator_0/4input_AND_0/not_0/in comparator_0/4input_AND_0/w_n8_2# 0.02fF
C1186 vdd comparator_0/4input_AND_2/w_68_n95# 0.02fF
C1187 AND_Block_0/and_1/a_n26_14# b1out_3 0.31fF
C1188 AND_Block_0/and_0/a_n26_14# AND_Block_0/and_0/w_26_9# 0.09fF
C1189 comparator_0/not_1/w_n2_10# b1out_2 0.09fF
C1190 4bitadder_0/fulladder_1/XOR_0/w_62_n20# 4bitadder_0/fulladder_1/axorb 0.04fF
C1191 comparator_0/a2xnorb2 gnd 1.27fF
C1192 comparator_0/4input_AND_2/w_n47_52# comparator_0/a3xnorb3 0.04fF
C1193 comparator_0/3input_AND_0/w_n14_24# comparator_0/b2bar 0.16fF
C1194 b3 enable_2/and_7/a_n26_14# 0.31fF
C1195 enable_2/a2 enable_2/and_2/a_n26_14# 0.31fF
C1196 4bitadder_1/fulladder_2/axorb 4bitadder_1/fulladder_2/XOR_1/w_62_37# 0.02fF
C1197 4bitadder_1/c2 4bitadder_1/fulladder_2/XOR_1/w_16_n1# 0.11fF
C1198 comparator_0/5input_AND_0/w_68_n82# comparator_0/a2xnorb2 0.16fF
C1199 a1out_1 4bitadder_1/fulladder_1/XOR_0/abar 0.13fF
C1200 enable_1/and_5/a_n26_14# enable_1/and_5/w_26_9# 0.09fF
C1201 enable_2/and_1/w_n43_8# enable_2/and_1/a_n26_14# 0.02fF
C1202 enable_1/and_2/a_n26_14# a2 0.31fF
C1203 enable_3/and_3/w_n43_8# enable_3/and_3/a_n26_14# 0.02fF
C1204 4bitadder_1/b0xorM 4bitadder_1/XOR_0/w_62_37# 0.02fF
C1205 4bitadder_1/c2 4bitadder_1/fulladder_2/XOR_1/abar 0.27fF
C1206 b2out_0 vdd 0.05fF
C1207 comparator_0/4input_OR_0/NOT_0/w_n2_10# vdd 0.18fF
C1208 4bitadder_0/fulladder_3/and_0/w_n43_8# vdd 0.07fF
C1209 4bitadder_0/fulladder_3/or_0/a_n15_32# 4bitadder_0/fulladder_3/or_0/w_58_101# 0.13fF
C1210 4bitadder_0/c2 4bitadder_0/fulladder_2/XOR_1/w_16_n1# 0.11fF
C1211 vdd 4bitadder_1/fulladder_3/and_1/w_n43_8# 0.07fF
C1212 enable_3/and_4/w_26_9# vdd 0.03fF
C1213 4bitadder_1/fulladder_2/or_0/w_58_101# 4bitadder_1/c3 0.02fF
C1214 enable_3/and_0/w_n43_8# vdd 0.07fF
C1215 comparator_0/b0bar comparator_0/a2xnorb2 0.38fF
C1216 s1 decoder_0/and_3/a_n26_14# 0.31fF
C1217 vdd 4bitadder_1/fulladder_2/or_0/a 0.14fF
C1218 comparator_0/4input_OR_0/w_n58_n43# comparator_0/t8 0.13fF
C1219 4bitadder_0/c2 4bitadder_0/fulladder_2/XOR_1/abar 0.27fF
C1220 4bitadder_1/fulladder_3/and_0/w_26_9# 4bitadder_1/fulladder_3/or_0/a 0.03fF
C1221 4bitadder_1/fulladder_0/or_0/w_n48_101# 4bitadder_1/fulladder_0/or_0/a 0.12fF
C1222 gnd decoder_0/and_1/b 0.19fF
C1223 4bitadder_0/b0xorM gnd 0.42fF
C1224 enable_2/and_0/w_n43_8# enable_2/en 0.09fF
C1225 4bitadder_0/fulladder_1/or_0/w_n48_101# 4bitadder_0/fulladder_1/or_0/a 0.12fF
C1226 4bitadder_0/fulladder_1/XOR_0/abar gnd 0.15fF
C1227 s0 4bitadder_1/XOR_2/w_16_n1# 0.11fF
C1228 a2out_2 comparator_0/a3xnorb3 0.60fF
C1229 comparator_0/xnor_0/not_0/w_n2_10# comparator_0/a3xnorb3 0.03fF
C1230 4bitadder_0/XOR_1/out s0 0.15fF
C1231 4bitadder_1/fulladder_2/and_1/w_26_9# 4bitadder_1/fulladder_2/and_1/a_n26_14# 0.09fF
C1232 4bitadder_0/fulladder_0/XOR_0/w_62_37# a0out_0 0.02fF
C1233 4bitadder_0/fulladder_0/and_0/w_n43_8# vdd 0.07fF
C1234 b2out_2 b1out_2 0.42fF
C1235 enable_1/and_1/w_26_9# vdd 0.03fF
C1236 s0 4bitadder_1/XOR_2/abar 0.28fF
C1237 a2out_2 comparator_0/a1xnorb1 0.46fF
C1238 4bitadder_0/fulladder_1/XOR_0/w_62_n20# 4bitadder_0/fulladder_1/XOR_0/abar 0.02fF
C1239 boout_2 comparator_0/xnor_3/XOR_0/bbar 0.02fF
C1240 4bitadder_1/XOR_1/w_n34_n1# 4bitadder_1/XOR_1/abar 0.03fF
C1241 4bitadder_1/XOR_0/abar s0 1.07fF
C1242 gnd 4bitadder_1/c3 0.91fF
C1243 AND_Block_0/and_3/w_26_9# vdd 0.03fF
C1244 b3 a3 0.31fF
C1245 vdd 4bitadder_1/fulladder_3/axorb 0.15fF
C1246 vdd comparator_0/5input_AND_1/w_31_n55# 0.06fF
C1247 a2out_1 b3out_1 0.33fF
C1248 s2_add vdd 0.19fF
C1249 4bitadder_0/XOR_1/w_n34_n1# 4bitadder_0/XOR_1/abar 0.03fF
C1250 4bitadder_1/fulladder_0/and_0/w_n43_8# s0 0.09fF
C1251 4bitadder_0/c3 4bitadder_0/fulladder_3/axorb 0.60fF
C1252 4bitadder_0/fulladder_2/and_1/w_n43_8# 4bitadder_0/XOR_2/out 0.09fF
C1253 4bitadder_1/fulladder_3/or_0/a_n15_32# 4bitadder_1/fulladder_3/or_0/w_58_101# 0.13fF
C1254 4bitadder_1/XOR_3/w_n34_n1# 4bitadder_1/XOR_3/abar 0.03fF
C1255 4bitadder_1/XOR_3/w_16_n1# 4bitadder_1/XOR_3/bbar 0.03fF
C1256 comparator_0/4input_OR_0/y comparator_0/t6 0.18fF
C1257 enable_0/and_6/w_n43_8# b2 0.09fF
C1258 4bitadder_0/XOR_2/w_n34_n1# vdd 0.02fF
C1259 vdd comparator_0/and_0/w_26_9# 0.03fF
C1260 4bitadder_0/XOR_3/w_n34_n1# 4bitadder_0/XOR_3/abar 0.03fF
C1261 4bitadder_0/XOR_3/w_16_n1# 4bitadder_0/XOR_3/bbar 0.03fF
C1262 enable_0/en gnd 0.01fF
C1263 s3_add vdd 0.10fF
C1264 4bitadder_0/fulladder_3/or_0/a_n15_32# 4bitadder_0/fulladder_3/or_0/w_n48_101# 0.05fF
C1265 enable_1/and_2/w_26_9# enable_1/and_2/a_n26_14# 0.09fF
C1266 a1out_1 a0_out1 1.88fF
C1267 vdd comparator_0/4input_AND_0/w_n47_52# 0.02fF
C1268 4bitadder_0/fulladder_2/XOR_0/w_62_37# 4bitadder_0/XOR_2/out 0.13fF
C1269 4bitadder_0/XOR_3/w_62_37# s0 0.13fF
C1270 vdd decoder_0/not_1/w_n2_10# 0.18fF
C1271 vdd 4bitadder_1/fulladder_3/XOR_0/w_n34_n1# 0.02fF
C1272 enable_3/and_3/w_n43_8# vdd 0.07fF
C1273 4bitadder_1/fulladder_3/and_1/w_n43_8# 4bitadder_1/XOR_3/out 0.09fF
C1274 b2out_0 s0 0.30fF
C1275 a3out_2 a0out_2 0.60fF
C1276 b2out_3 gnd 0.24fF
C1277 enable_1/and_3/a_n26_14# a3 0.31fF
C1278 b0out_0 4bitadder_0/XOR_0/abar 0.13fF
C1279 4bitadder_0/fulladder_3/and_1/w_n43_8# 4bitadder_0/XOR_3/out 0.09fF
C1280 enable_3/and_4/w_n43_8# enable_3/and_4/a_n26_14# 0.02fF
C1281 comparator_0/4input_AND_1/not_0/in comparator_0/4input_AND_1/w_n8_2# 0.02fF
C1282 b2out_3 AND_Block_0/and_2/w_n43_8# 0.09fF
C1283 a1 enable_2/en 0.28fF
C1284 enable_1/and_7/w_26_9# enable_1/and_7/a_n26_14# 0.09fF
C1285 4bitadder_0/fulladder_3/axorb 4bitadder_0/fulladder_3/XOR_1/abar 0.13fF
C1286 comparator_0/a1xnorb1 comparator_0/4input_AND_0/not_0/in 0.18fF
C1287 comparator_0/4input_AND_1/not_0/in comparator_0/a3xnorb3 0.18fF
C1288 enable_2/en enable_2/and_3/w_n43_8# 0.09fF
C1289 b2 enable_2/and_6/w_n43_8# 0.09fF
C1290 a2out_2 b2out_2 0.46fF
C1291 vdd comparator_0/4input_AND_1/not_0/w_n2_10# 0.18fF
C1292 comparator_0/xnor_1/XOR_0/w_n34_n1# comparator_0/xnor_1/XOR_0/abar 0.03fF
C1293 comparator_0/xnor_1/XOR_0/w_16_n1# comparator_0/xnor_1/XOR_0/bbar 0.03fF
C1294 comparator_0/xnor_1/XOR_0/w_62_n20# comparator_0/xnor_1/not_0/in 0.04fF
C1295 comparator_0/4input_OR_0/y comparator_0/4input_OR_0/w_n58_n43# 0.02fF
C1296 4bitadder_0/fulladder_2/axorb 4bitadder_0/c2 0.54fF
C1297 enable_2/and_6/a_n26_14# enable_2/and_6/w_n43_8# 0.02fF
C1298 4bitadder_0/fulladder_0/and_1/w_26_9# 4bitadder_0/fulladder_0/and_1/a_n26_14# 0.09fF
C1299 4bitadder_1/XOR_0/w_62_n20# 4bitadder_1/XOR_0/abar 0.02fF
C1300 vdd a2out_1 0.33fF
C1301 AND_Block_0/and_3/w_n43_8# b3out_3 0.09fF
C1302 boout_2 gnd 0.90fF
C1303 4bitadder_0/fulladder_1/or_0/a_n15_32# 4bitadder_0/fulladder_1/or_0/b 0.19fF
C1304 enable_2/and_6/a_n26_14# enable_2/and_6/w_26_9# 0.09fF
C1305 4bitadder_0/XOR_0/w_62_n20# 4bitadder_0/XOR_0/abar 0.02fF
C1306 4bitadder_0/fulladder_1/XOR_1/w_16_n1# vdd 0.02fF
C1307 gnd b3out_1 0.62fF
C1308 b1 gnd 0.21fF
C1309 a2out_0 gnd 1.02fF
C1310 comparator_0/t4 comparator_0/t1 0.18fF
C1311 a2out_1 b0out_1 0.09fF
C1312 4bitadder_1/fulladder_3/axorb 4bitadder_1/XOR_3/out 0.13fF
C1313 4bitadder_0/fulladder_0/and_0/w_n43_8# s0 0.09fF
C1314 vdd 4bitadder_1/fulladder_1/XOR_1/w_16_n1# 0.02fF
C1315 4bitadder_1/fulladder_1/XOR_0/w_n34_n1# a1out_1 0.11fF
C1316 4bitadder_0/fulladder_1/or_0/a_n15_32# 4bitadder_0/fulladder_1/or_0/w_58_101# 0.13fF
C1317 4bitadder_0/fulladder_0/axorb 4bitadder_0/fulladder_0/and_0/w_n43_8# 0.09fF
C1318 comparator_0/4input_OR_1/y comparator_0/t1 0.18fF
C1319 4bitadder_1/XOR_1/out 4bitadder_1/fulladder_1/XOR_0/w_62_37# 0.13fF
C1320 enable_3/and_5/w_26_9# vdd 0.03fF
C1321 4bitadder_1/fulladder_2/axorb 4bitadder_1/fulladder_2/XOR_0/w_62_37# 0.02fF
C1322 4bitadder_0/fulladder_2/or_0/w_58_101# vdd 0.05fF
C1323 a1out_2 comparator_0/not_5/w_n2_10# 0.09fF
C1324 comparator_0/xnor_3/XOR_0/w_n34_n1# comparator_0/xnor_3/XOR_0/abar 0.03fF
C1325 4bitadder_0/fulladder_2/XOR_0/bbar 4bitadder_0/XOR_2/out 0.02fF
C1326 4bitadder_0/fulladder_1/and_0/w_n43_8# 4bitadder_0/c1 0.09fF
C1327 a3out_0 gnd 0.99fF
C1328 enable_3/and_7/w_n43_8# enable_3/and_7/a_n26_14# 0.02fF
C1329 vdd 4bitadder_1/fulladder_2/or_0/w_58_101# 0.05fF
C1330 comparator_0/t1 comparator_0/t3 0.18fF
C1331 4bitadder_0/fulladder_1/axorb 4bitadder_0/fulladder_1/XOR_1/w_62_37# 0.02fF
C1332 b3out_0 4bitadder_0/XOR_3/abar 0.13fF
C1333 4bitadder_1/fulladder_0/axorb 4bitadder_1/fulladder_0/XOR_1/w_62_37# 0.02fF
C1334 4bitadder_1/c1 4bitadder_1/fulladder_1/XOR_1/bbar 0.02fF
C1335 vdd comparator_0/xnor_0/XOR_0/w_16_n1# 0.02fF
C1336 4bitadder_1/fulladder_3/XOR_0/w_62_37# a3out_1 0.02fF
C1337 boout_2 comparator_0/a2xnorb2 0.69fF
C1338 enable_0/and_1/w_26_9# vdd 0.03fF
C1339 4bitadder_1/fulladder_2/or_0/w_n48_101# 4bitadder_1/fulladder_2/or_0/b 0.12fF
C1340 4bitadder_0/fulladder_2/XOR_1/w_n34_n1# 4bitadder_0/fulladder_2/XOR_1/abar 0.03fF
C1341 4bitadder_0/fulladder_2/XOR_1/w_16_n1# 4bitadder_0/fulladder_2/XOR_1/bbar 0.03fF
C1342 4bitadder_0/fulladder_2/XOR_1/w_62_n20# s2_add 0.04fF
C1343 AND_Block_0/and_3/w_n43_8# a3out_3 0.09fF
C1344 enable_2/and_2/w_26_9# a2out_2 0.03fF
C1345 4bitadder_1/fulladder_3/axorb 4bitadder_1/fulladder_3/and_0/w_n43_8# 0.09fF
C1346 a2 gnd 0.21fF
C1347 comparator_0/xnor_0/not_0/in gnd 0.03fF
C1348 4bitadder_0/XOR_2/bbar s0 0.02fF
C1349 4bitadder_0/c3 4bitadder_0/fulladder_3/XOR_1/bbar 0.02fF
C1350 4bitadder_0/fulladder_3/XOR_0/w_62_37# a3out_0 0.02fF
C1351 enable_1/and_3/w_26_9# enable_1/and_3/a_n26_14# 0.09fF
C1352 4bitadder_1/fulladder_0/XOR_0/abar 4bitadder_1/b0xorM 0.25fF
C1353 comparator_0/5input_AND_0/not_0/in comparator_0/5input_AND_0/w_n37_15# 0.05fF
C1354 4bitadder_1/fulladder_3/XOR_0/bbar 4bitadder_1/XOR_3/out 0.02fF
C1355 4bitadder_0/fulladder_0/or_0/w_58_101# vdd 0.05fF
C1356 enable_1/and_2/w_26_9# a2out_1 0.03fF
C1357 4bitadder_0/fulladder_3/XOR_0/bbar 4bitadder_0/XOR_3/out 0.02fF
C1358 vdd gnd 5.30fF
C1359 enable_1/and_1/w_n43_8# vdd 0.07fF
C1360 vdd comparator_0/5input_AND_0/w_68_n82# 0.05fF
C1361 vdd comparator_0/not_3/w_n2_10# 0.18fF
C1362 enable_1/and_4/a_n26_14# b0 0.31fF
C1363 a0 a1 0.31fF
C1364 vdd comparator_0/4input_AND_1/w_n47_52# 0.02fF
C1365 AND_Block_0/and_2/w_n43_8# vdd 0.07fF
C1366 comparator_0/b3 comparator_0/a1xnorb1 0.42fF
C1367 AND_Block_0/and_1/w_26_9# out1 0.03fF
C1368 a3 enable_2/en 0.28fF
C1369 4bitadder_0/fulladder_1/and_1/w_26_9# vdd 0.03fF
C1370 4bitadder_1/fulladder_3/XOR_1/w_n34_n1# 4bitadder_1/fulladder_3/XOR_1/abar 0.03fF
C1371 4bitadder_1/fulladder_3/XOR_1/w_16_n1# 4bitadder_1/fulladder_3/XOR_1/bbar 0.03fF
C1372 4bitadder_1/fulladder_3/XOR_1/w_62_n20# s3_sub 0.04fF
C1373 vdd 4bitadder_1/fulladder_0/and_0/w_26_9# 0.03fF
C1374 enable_1/and_6/w_n43_8# vdd 0.07fF
C1375 a1out_3 gnd 0.18fF
C1376 a2out_1 s0 0.22fF
C1377 AND_Block_0/and_2/w_26_9# vdd 0.03fF
C1378 gnd b0out_1 0.14fF
C1379 4bitadder_1/XOR_2/w_n34_n1# b2out_1 0.11fF
C1380 4bitadder_0/fulladder_1/or_0/b gnd 0.37fF
C1381 enable_1/en gnd 0.13fF
C1382 4bitadder_1/fulladder_0/and_1/w_n43_8# a0_out1 0.09fF
C1383 4bitadder_0/fulladder_3/XOR_1/w_n34_n1# 4bitadder_0/fulladder_3/XOR_1/abar 0.03fF
C1384 4bitadder_0/fulladder_3/XOR_1/w_16_n1# 4bitadder_0/fulladder_3/XOR_1/bbar 0.03fF
C1385 4bitadder_0/fulladder_3/XOR_1/w_62_n20# s3_add 0.04fF
C1386 4bitadder_0/fulladder_0/XOR_1/abar gnd 0.15fF
C1387 AND_Block_0/and_0/w_n43_8# AND_Block_0/and_0/a_n26_14# 0.02fF
C1388 enable_1/and_1/w_n43_8# enable_1/en 0.09fF
C1389 vdd comparator_0/4input_OR_1/w_n58_n43# 0.03fF
C1390 comparator_0/xnor_2/XOR_0/w_n34_n1# a1out_2 0.11fF
C1391 4bitadder_0/fulladder_2/or_0/w_n48_101# vdd 0.05fF
C1392 enable_1/and_6/w_26_9# vdd 0.03fF
C1393 vdd comparator_0/5input_AND_1/not_0/w_n2_10# 0.17fF
C1394 gnd 4bitadder_1/fulladder_1/or_0/b 0.37fF
C1395 a1out_2 comparator_0/a3xnorb3 0.53fF
C1396 comparator_0/b0bar comparator_0/5input_AND_0/w_n4_n20# 0.18fF
C1397 4bitadder_0/XOR_1/out a1out_0 1.87fF
C1398 4bitadder_0/fulladder_1/and_1/w_26_9# 4bitadder_0/fulladder_1/or_0/b 0.03fF
C1399 enable_0/and_7/w_26_9# vdd 0.03fF
C1400 vdd comparator_0/b0bar 0.14fF
C1401 4bitadder_1/XOR_2/w_62_n20# 4bitadder_1/XOR_2/abar 0.02fF
C1402 vdd 4bitadder_1/XOR_0/w_16_n1# 0.02fF
C1403 vdd comparator_0/and_1/w_n43_8# 0.07fF
C1404 enable_1/and_6/w_n43_8# enable_1/en 0.09fF
C1405 enable_1/and_5/w_n43_8# enable_1/and_5/a_n26_14# 0.02fF
C1406 b2 b3 0.33fF
C1407 AND_Block_0/and_0/a_n26_14# b0out_3 0.31fF
C1408 vdd 4bitadder_1/fulladder_0/or_0/w_58_101# 0.05fF
C1409 vdd decoder_0/and_3/w_26_9# 0.03fF
C1410 comparator_0/xnor_2/XOR_0/w_62_n20# comparator_0/xnor_2/XOR_0/abar 0.02fF
C1411 4bitadder_0/fulladder_1/axorb vdd 0.15fF
C1412 enable_0/and_3/w_26_9# a3out_0 0.03fF
C1413 4bitadder_0/XOR_2/w_62_n20# 4bitadder_0/XOR_2/abar 0.02fF
C1414 comparator_0/a1xnorb1 a1out_2 0.54fF
C1415 4bitadder_0/fulladder_2/and_0/w_n43_8# 4bitadder_0/fulladder_2/and_0/a_n26_14# 0.02fF
C1416 enable_0/en enable_0/and_2/w_n43_8# 0.09fF
C1417 enable_0/and_1/w_n43_8# a1 0.09fF
C1418 vdd comparator_0/4input_AND_2/w_n8_2# 0.02fF
C1419 4bitadder_1/XOR_1/out gnd 0.42fF
C1420 4bitadder_0/c3 4bitadder_0/fulladder_3/and_0/a_n26_14# 0.10fF
C1421 4bitadder_1/XOR_0/abar 4bitadder_1/XOR_0/w_n34_n1# 0.03fF
C1422 4bitadder_1/fulladder_1/and_1/w_n43_8# 4bitadder_1/fulladder_1/and_1/a_n26_14# 0.02fF
C1423 4bitadder_0/fulladder_0/XOR_0/w_16_n1# 4bitadder_0/b0xorM 0.11fF
C1424 vdd decoder_0/not_0/w_n2_10# 0.18fF
C1425 4bitadder_1/c2 4bitadder_1/fulladder_2/XOR_1/w_62_37# 0.13fF
C1426 a1out_1 4bitadder_1/fulladder_1/and_1/w_n43_8# 0.09fF
C1427 comparator_0/a0xnorb0 comparator_0/a3xnorb3 0.29fF
C1428 vdd comparator_0/a2xnorb2 2.46fF
C1429 b0out_3 b1out_3 24.79fF
C1430 4bitadder_0/XOR_0/abar 4bitadder_0/XOR_0/w_n34_n1# 0.03fF
C1431 4bitadder_1/fulladder_1/and_0/a_n26_14# 4bitadder_1/fulladder_1/and_0/w_n43_8# 0.02fF
C1432 4bitadder_0/XOR_1/out 4bitadder_0/XOR_1/w_62_n20# 0.04fF
C1433 b3 enable_2/b1 0.13fF
C1434 4bitadder_0/XOR_1/abar s0 0.25fF
C1435 4bitadder_1/c2 s2_sub 0.04fF
C1436 comparator_0/a1xnorb1 comparator_0/a0xnorb0 0.40fF
C1437 a2out_1 b1out_1 0.12fF
C1438 4bitadder_1/fulladder_3/XOR_0/w_62_n20# 4bitadder_1/fulladder_3/XOR_0/abar 0.02fF
C1439 comparator_0/4input_AND_2/not_0/w_n2_10# comparator_0/t3 0.03fF
C1440 4bitadder_0/fulladder_2/axorb 4bitadder_0/fulladder_2/XOR_1/w_n34_n1# 0.11fF
C1441 4bitadder_0/c2 4bitadder_0/fulladder_2/XOR_1/w_62_37# 0.13fF
C1442 enable_2/and_3/w_26_9# vdd 0.03fF
C1443 comparator_0/b3 b2out_2 0.43fF
C1444 comparator_0/t2 comparator_0/3input_AND_1/not_0/w_n2_10# 0.03fF
C1445 4bitadder_0/XOR_2/out 4bitadder_0/XOR_2/w_62_37# 0.02fF
C1446 4bitadder_0/fulladder_3/XOR_0/w_62_n20# 4bitadder_0/fulladder_3/XOR_0/abar 0.02fF
C1447 enable_0/and_3/w_26_9# vdd 0.03fF
C1448 comparator_0/4input_AND_2/not_0/in comparator_0/4input_AND_2/w_68_n95# 0.02fF
C1449 comparator_0/b3bar comparator_0/and_0/a_n26_14# 0.10fF
C1450 enable_1/and_6/a_n26_14# b2 0.31fF
C1451 enable_0/en b1 0.34fF
C1452 gnd 4bitadder_1/XOR_3/out 0.42fF
C1453 4bitadder_0/c2 s2_add 0.04fF
C1454 enable_1/and_4/w_26_9# enable_1/and_4/a_n26_14# 0.09fF
C1455 b0 gnd 0.30fF
C1456 4bitadder_1/fulladder_1/or_0/w_n48_101# 4bitadder_1/fulladder_1/or_0/a 0.12fF
C1457 comparator_0/xnor_1/not_0/w_n2_10# comparator_0/xnor_1/not_0/in 0.09fF
C1458 vdd 4bitadder_1/fulladder_1/and_0/w_26_9# 0.03fF
C1459 vdd decoder_0/and_1/b 0.04fF
C1460 comparator_0/t1 comparator_0/t2 0.18fF
C1461 gnd s0 8.09fF
C1462 s0 4bitadder_1/XOR_2/w_62_37# 0.13fF
C1463 4bitadder_0/fulladder_0/axorb gnd 0.09fF
C1464 4bitadder_0/fulladder_3/and_0/w_n43_8# 4bitadder_0/fulladder_3/axorb 0.09fF
C1465 vdd comparator_0/4input_OR_1/NOT_0/w_n2_10# 0.18fF
C1466 4bitadder_1/fulladder_2/and_1/w_n43_8# a2out_1 0.09fF
C1467 a0 a3 0.31fF
C1468 enable_1/and_0/w_26_9# a0_out1 0.03fF
C1469 a2out_2 b1out_2 1.07fF
C1470 b2out_2 a1out_2 0.65fF
C1471 4bitadder_0/fulladder_2/XOR_0/w_n34_n1# a2out_0 0.11fF
C1472 4bitadder_0/fulladder_1/and_0/w_26_9# vdd 0.03fF
C1473 enable_2/a0 gnd 0.07fF
C1474 comparator_0/xnor_3/XOR_0/w_62_n20# comparator_0/xnor_3/XOR_0/abar 0.02fF
C1475 b3 enable_2/a2 0.10fF
C1476 vdd 4bitadder_1/c3 0.12fF
C1477 4bitadder_1/fulladder_0/XOR_1/abar s0 0.27fF
C1478 vdd comparator_0/5input_AND_1/w_n37_15# 0.05fF
C1479 4bitadder_0/fulladder_0/XOR_0/w_n34_n1# a0out_0 0.11fF
C1480 enable_1/and_7/w_n43_8# vdd 0.07fF
C1481 comparator_0/4input_OR_1/NOT_0/w_n2_10# bga 0.03fF
C1482 enable_1/and_0/a_n26_14# enable_1/and_0/w_n43_8# 0.02fF
C1483 enable_3/and_5/w_n43_8# b1 0.09fF
C1484 4bitadder_1/XOR_0/w_16_n1# s0 0.11fF
C1485 4bitadder_1/fulladder_1/axorb 4bitadder_1/fulladder_1/XOR_1/w_n34_n1# 0.11fF
C1486 comparator_0/b1bar comparator_0/4input_AND_1/not_0/in 0.18fF
C1487 a3out_2 comparator_0/and_0/w_n43_8# 0.09fF
C1488 comparator_0/5input_AND_1/not_0/in comparator_0/5input_AND_1/w_68_n82# 0.02fF
C1489 4bitadder_1/fulladder_3/and_0/a_n26_14# 4bitadder_1/c3 0.10fF
C1490 4bitadder_0/fulladder_1/XOR_1/w_62_37# s1_add 0.02fF
C1491 enable_0/and_6/w_26_9# enable_0/and_6/a_n26_14# 0.09fF
C1492 4bitadder_1/fulladder_3/axorb 4bitadder_1/fulladder_3/XOR_1/abar 0.13fF
C1493 4bitadder_0/XOR_1/w_62_37# s0 0.13fF
C1494 4bitadder_0/fulladder_3/and_0/w_26_9# vdd 0.03fF
C1495 enable_0/en a2 0.38fF
C1496 enable_3/and_7/w_26_9# b3out_3 0.03fF
C1497 comparator_0/not_7/w_n2_10# comparator_0/a3bar 0.03fF
C1498 4bitadder_1/fulladder_2/or_0/w_n48_101# 4bitadder_1/fulladder_2/or_0/a 0.12fF
C1499 comparator_0/5input_AND_1/w_106_n113# comparator_0/a3xnorb3 0.17fF
C1500 enable_1/and_7/w_n43_8# enable_1/en 0.09fF
C1501 enable_2/and_5/w_26_9# b1out_2 0.03fF
C1502 enable_0/en enable_0/and_4/w_n43_8# 0.09fF
C1503 enable_0/and_2/w_n43_8# a2 0.09fF
C1504 s0 decoder_0/not_0/w_n2_10# 0.09fF
C1505 gnd b1out_1 1.08fF
C1506 enable_3/en b3 0.32fF
C1507 enable_0/en vdd 0.93fF
C1508 enable_0/and_6/a_n26_14# b2 0.31fF
C1509 4bitadder_1/fulladder_1/XOR_1/w_62_37# s1_sub 0.02fF
C1510 vdd equal 0.04fF
C1511 4bitadder_0/fulladder_2/XOR_0/w_16_n1# 4bitadder_0/XOR_2/out 0.11fF
C1512 enable_2/and_2/w_n43_8# vdd 0.07fF
C1513 4bitadder_0/XOR_1/w_n34_n1# vdd 0.02fF
C1514 AND_Block_0/and_1/w_n43_8# b1out_3 0.09fF
C1515 a2out_0 a3out_0 1.82fF
C1516 vdd comparator_0/3input_AND_0/w_32_n21# 0.03fF
C1517 4bitadder_0/fulladder_3/axorb 4bitadder_0/fulladder_3/XOR_1/w_62_37# 0.02fF
C1518 enable_0/and_2/w_n43_8# vdd 0.07fF
C1519 enable_2/and_7/w_n43_8# b3 0.09fF
C1520 4bitadder_0/fulladder_3/or_0/a_n15_32# 4bitadder_0/fulladder_3/or_0/b 0.19fF
C1521 b2out_3 vdd 0.14fF
C1522 comparator_0/3input_AND_1/not_0/in comparator_0/3input_AND_1/w_69_n71# 0.02fF
C1523 4bitadder_0/fulladder_2/XOR_0/w_n34_n1# vdd 0.02fF
C1524 enable_3/en enable_3/and_2/w_n43_8# 0.09fF
C1525 4bitadder_1/fulladder_0/axorb 4bitadder_1/b0xorM 0.13fF
C1526 4bitadder_1/fulladder_0/XOR_1/w_62_n20# 4bitadder_1/fulladder_0/XOR_1/abar 0.02fF
C1527 comparator_0/xnor_1/XOR_0/w_16_n1# b2out_2 0.11fF
C1528 4bitadder_0/fulladder_2/XOR_0/w_62_37# 4bitadder_0/fulladder_2/axorb 0.02fF
C1529 4bitadder_0/fulladder_0/XOR_0/abar gnd 0.15fF
C1530 4bitadder_0/fulladder_0/and_1/w_n43_8# a0out_0 0.09fF
C1531 4bitadder_1/fulladder_2/XOR_0/w_n34_n1# a2out_1 0.11fF
C1532 4bitadder_1/fulladder_2/XOR_0/w_16_n1# 4bitadder_1/XOR_2/out 0.11fF
C1533 a0out_2 gnd 0.56fF
C1534 b1 a2 0.19fF
C1535 s0 decoder_0/and_1/b 0.19fF
C1536 comparator_0/a1xnorb1 comparator_0/4input_AND_0/w_29_n46# 0.16fF
C1537 4bitadder_0/b0xorM s0 0.26fF
C1538 b2 enable_2/en 0.29fF
C1539 enable_2/and_0/a_n26_14# enable_2/a0 0.31fF
C1540 vdd boout_2 0.94fF
C1541 comparator_0/and_0/w_n43_8# comparator_0/b3bar 0.09fF
C1542 comparator_0/and_0/w_26_9# comparator_0/and_0/a_n26_14# 0.09fF
C1543 enable_3/and_5/w_n43_8# vdd 0.07fF
C1544 b2out_2 comparator_0/xnor_1/XOR_0/abar 0.30fF
C1545 s0 4bitadder_1/XOR_1/bbar 0.02fF
C1546 4bitadder_0/fulladder_0/axorb 4bitadder_0/b0xorM 0.13fF
C1547 4bitadder_1/fulladder_2/XOR_0/abar 4bitadder_1/XOR_2/out 0.25fF
C1548 vdd b3out_1 0.13fF
C1549 b1 vdd 0.35fF
C1550 decoder_0/not_1/w_n2_10# s1 0.09fF
C1551 4bitadder_1/c3 4bitadder_1/XOR_3/out 0.41fF
C1552 a2out_0 vdd 0.35fF
C1553 enable_2/and_5/w_n43_8# enable_2/en 0.09fF
C1554 s1_add vdd 0.19fF
C1555 gnd 4bitadder_1/XOR_3/abar 0.20fF
C1556 4bitadder_1/fulladder_1/axorb 4bitadder_1/c1 0.54fF
C1557 comparator_0/t5 comparator_0/t7 0.21fF
C1558 vdd 4bitadder_1/fulladder_0/XOR_0/w_n34_n1# 0.02fF
C1559 4bitadder_0/fulladder_2/or_0/a gnd 0.01fF
C1560 vdd enable_0/and_5/w_26_9# 0.03fF
C1561 vdd s1_sub 0.19fF
C1562 comparator_0/b0bar a0out_2 0.25fF
C1563 enable_2/en enable_2/b1 0.19fF
C1564 b3out_0 4bitadder_0/XOR_3/w_62_37# 0.02fF
C1565 4bitadder_1/fulladder_2/XOR_1/w_62_n20# 4bitadder_1/fulladder_2/XOR_1/bbar 0.13fF
C1566 comparator_0/xnor_3/XOR_0/w_62_37# boout_2 0.13fF
C1567 4bitadder_0/fulladder_2/XOR_0/w_62_n20# 4bitadder_0/fulladder_2/XOR_0/bbar 0.13fF
C1568 enable_1/en b1 0.25fF
C1569 comparator_0/xnor_0/XOR_0/w_62_37# comparator_0/xnor_0/not_0/in 0.02fF
C1570 a3out_0 vdd 0.29fF
C1571 gnd 4bitadder_1/fulladder_2/axorb 0.09fF
C1572 4bitadder_0/fulladder_0/XOR_0/w_16_n1# vdd 0.02fF
C1573 enable_0/and_1/w_n43_8# enable_0/and_1/a_n26_14# 0.02fF
C1574 4bitadder_1/fulladder_3/or_0/w_n48_101# 4bitadder_1/fulladder_3/or_0/a_n15_32# 0.05fF
C1575 agb vdd 0.04fF
C1576 4bitadder_0/c2 gnd 0.97fF
C1577 b2out_0 4bitadder_0/XOR_2/abar 0.13fF
C1578 a1 a3 0.31fF
C1579 comparator_0/b3 comparator_0/xnor_0/XOR_0/bbar 0.02fF
C1580 enable_0/en b0 0.38fF
C1581 4bitadder_0/fulladder_2/or_0/w_n48_101# 4bitadder_0/fulladder_2/or_0/a 0.12fF
C1582 a0out_2 comparator_0/a2xnorb2 0.38fF
C1583 a3 enable_2/and_3/w_n43_8# 0.09fF
C1584 enable_3/and_3/w_26_9# a3out_3 0.03fF
C1585 enable_3/and_1/w_n43_8# a1 0.09fF
C1586 4bitadder_1/c3 4bitadder_1/fulladder_3/and_0/w_n43_8# 0.09fF
C1587 comparator_0/b1bar a1out_2 0.18fF
C1588 enable_0/and_3/w_n43_8# a3 0.09fF
C1589 4bitadder_0/XOR_0/bbar s0 0.02fF
C1590 4bitadder_0/fulladder_0/or_0/a gnd 0.01fF
C1591 enable_3/and_0/a_n26_14# enable_3/and_0/w_n43_8# 0.02fF
C1592 a2 vdd 0.31fF
C1593 enable_2/and_4/w_n43_8# vdd 0.07fF
C1594 enable_0/and_1/w_26_9# a1out_0 0.03fF
C1595 a3out_2 comparator_0/a3xnorb3 0.18fF
C1596 enable_0/and_4/w_n43_8# vdd 0.07fF
C1597 vdd comparator_0/5input_AND_0/w_n4_n20# 0.05fF
C1598 enable_2/en enable_2/a2 0.17fF
C1599 comparator_0/b3 b1out_2 0.48fF
C1600 a3out_2 comparator_0/a1xnorb1 0.17fF
C1601 enable_0/and_4/w_26_9# b0out_0 0.03fF
C1602 comparator_0/a0bar comparator_0/a3xnorb3 0.29fF
C1603 enable_1/en a2 0.28fF
C1604 enable_1/and_1/w_26_9# enable_1/and_1/a_n26_14# 0.09fF
C1605 4bitadder_1/XOR_1/w_62_n20# 4bitadder_1/XOR_1/abar 0.02fF
C1606 vdd comparator_0/a2bar 0.45fF
C1607 4bitadder_0/fulladder_0/XOR_0/abar 4bitadder_0/b0xorM 0.25fF
C1608 4bitadder_0/fulladder_0/XOR_1/w_16_n1# vdd 0.02fF
C1609 enable_3/en enable_3/and_4/w_n43_8# 0.09fF
C1610 gnd 4bitadder_1/fulladder_3/XOR_1/abar 0.15fF
C1611 a1out_3 vdd 0.16fF
C1612 vdd 4bitadder_1/fulladder_1/or_0/w_58_101# 0.05fF
C1613 4bitadder_0/XOR_1/w_62_n20# 4bitadder_0/XOR_1/abar 0.02fF
C1614 a1out_0 gnd 0.92fF
C1615 vdd b0out_1 0.13fF
C1616 comparator_0/a0bar comparator_0/a1xnorb1 0.03fF
C1617 AND_Block_0/and_0/w_n43_8# a0out_3 0.09fF
C1618 b2 a0 0.31fF
C1619 a2out_3 b1out_3 0.12fF
C1620 comparator_0/5input_AND_1/not_0/in comparator_0/a3xnorb3 0.23fF
C1621 enable_2/and_0/a_n26_14# enable_2/and_0/w_26_9# 0.09fF
C1622 vdd 4bitadder_1/fulladder_0/and_1/w_26_9# 0.03fF
C1623 vdd bga 0.04fF
C1624 4bitadder_0/fulladder_3/and_0/a_n26_14# 4bitadder_0/fulladder_3/and_0/w_n43_8# 0.02fF
C1625 enable_1/en vdd 0.92fF
C1626 b1 b0 4.71fF
C1627 decoder_0/and_0/w_n43_8# decoder_0/and_0/a_n26_14# 0.02fF
C1628 a2out_2 comparator_0/not_6/w_n2_10# 0.09fF
C1629 comparator_0/4input_AND_1/w_29_n46# comparator_0/a3xnorb3 0.16fF
C1630 4bitadder_0/fulladder_3/axorb gnd 0.09fF
C1631 out2 gnd 0.01fF
C1632 4bitadder_0/fulladder_2/and_0/w_26_9# vdd 0.03fF
C1633 4bitadder_0/fulladder_1/and_1/w_n43_8# 4bitadder_0/fulladder_1/and_1/a_n26_14# 0.02fF
C1634 s0 b3out_1 0.19fF
C1635 4bitadder_1/XOR_2/w_n34_n1# 4bitadder_1/XOR_2/abar 0.03fF
C1636 4bitadder_1/XOR_2/w_16_n1# 4bitadder_1/XOR_2/bbar 0.03fF
C1637 gnd 4bitadder_1/fulladder_1/XOR_0/abar 0.15fF
C1638 a2out_0 s0 0.31fF
C1639 a0out_3 b0out_3 2.02fF
C1640 vdd decoder_0/and_2/w_n43_8# 0.07fF
C1641 comparator_0/a1xnorb1 comparator_0/5input_AND_1/not_0/in 0.23fF
C1642 4bitadder_0/fulladder_0/XOR_1/w_62_n20# 4bitadder_0/fulladder_0/XOR_1/bbar 0.13fF
C1643 4bitadder_0/fulladder_1/or_0/w_58_101# vdd 0.05fF
C1644 enable_3/and_7/w_n43_8# vdd 0.07fF
C1645 a1out_2 b1out_2 0.88fF
C1646 comparator_0/4input_AND_2/not_0/in gnd 0.24fF
C1647 comparator_0/xnor_2/XOR_0/w_n34_n1# comparator_0/xnor_2/XOR_0/abar 0.03fF
C1648 comparator_0/xnor_2/XOR_0/w_16_n1# comparator_0/xnor_2/XOR_0/bbar 0.03fF
C1649 comparator_0/xnor_2/XOR_0/w_62_n20# comparator_0/xnor_2/not_0/in 0.04fF
C1650 4bitadder_0/XOR_2/w_n34_n1# 4bitadder_0/XOR_2/abar 0.03fF
C1651 4bitadder_0/XOR_2/w_16_n1# 4bitadder_0/XOR_2/bbar 0.03fF
C1652 enable_3/and_7/w_26_9# enable_3/and_7/a_n26_14# 0.09fF
C1653 gnd s1 0.34fF
C1654 comparator_0/and_0/a_n26_14# gnd 0.00fF
C1655 AND_Block_0/and_2/w_26_9# out2 0.03fF
C1656 a1 enable_2/and_1/a_n26_14# 0.31fF
C1657 4bitadder_1/fulladder_3/or_0/w_n48_101# 4bitadder_1/fulladder_3/or_0/b 0.12fF
C1658 comparator_0/3input_AND_0/not_0/in gnd 0.21fF
C1659 enable_2/and_7/w_n43_8# enable_2/en 0.09fF
C1660 4bitadder_1/fulladder_0/XOR_1/w_n34_n1# 4bitadder_1/fulladder_0/XOR_1/abar 0.03fF
C1661 comparator_0/xnor_1/not_0/w_n2_10# comparator_0/a2xnorb2 0.03fF
C1662 enable_2/and_2/w_n43_8# enable_2/and_2/a_n26_14# 0.02fF
C1663 a3out_0 s0 0.08fF
C1664 vdd comparator_0/t6 0.04fF
C1665 enable_0/and_1/a_n26_14# a1 0.31fF
C1666 4bitadder_0/c1 4bitadder_0/XOR_1/out 0.37fF
C1667 4bitadder_0/fulladder_3/axorb 4bitadder_0/fulladder_3/XOR_0/w_62_37# 0.02fF
C1668 enable_0/and_5/a_n26_14# b1 0.31fF
C1669 decoder_0/and_3/a_n26_14# Gnd 0.05fF
C1670 s1 Gnd 1.48fF
C1671 decoder_0/and_3/w_26_9# Gnd 0.82fF
C1672 decoder_0/and_3/w_n43_8# Gnd 0.82fF
C1673 decoder_0/and_2/a_n26_14# Gnd 0.05fF
C1674 decoder_0/and_2/w_26_9# Gnd 0.82fF
C1675 decoder_0/and_2/w_n43_8# Gnd 0.82fF
C1676 decoder_0/and_1/a_n26_14# Gnd 0.05fF
C1677 decoder_0/and_1/w_26_9# Gnd 0.82fF
C1678 decoder_0/and_1/w_n43_8# Gnd 0.82fF
C1679 decoder_0/and_0/a_n26_14# Gnd 0.05fF
C1680 decoder_0/and_0/w_26_9# Gnd 0.82fF
C1681 decoder_0/and_0/w_n43_8# Gnd 0.82fF
C1682 decoder_0/not_1/w_n2_10# Gnd 0.90fF
C1683 decoder_0/not_0/w_n2_10# Gnd 0.90fF
C1684 4bitadder_1/XOR_3/abar Gnd 0.11fF
C1685 4bitadder_1/XOR_3/bbar Gnd 0.06fF
C1686 4bitadder_1/XOR_3/w_62_n20# Gnd 0.87fF
C1687 4bitadder_1/XOR_3/w_16_n1# Gnd 0.75fF
C1688 4bitadder_1/XOR_3/w_n34_n1# Gnd 0.75fF
C1689 4bitadder_1/XOR_3/w_62_37# Gnd 0.72fF
C1690 4bitadder_1/XOR_2/abar Gnd 0.11fF
C1691 4bitadder_1/XOR_2/bbar Gnd 0.06fF
C1692 4bitadder_1/XOR_2/w_62_n20# Gnd 0.87fF
C1693 4bitadder_1/XOR_2/w_16_n1# Gnd 0.75fF
C1694 4bitadder_1/XOR_2/w_n34_n1# Gnd 0.75fF
C1695 4bitadder_1/XOR_2/w_62_37# Gnd 0.72fF
C1696 4bitadder_1/XOR_1/abar Gnd 0.11fF
C1697 4bitadder_1/XOR_1/bbar Gnd 0.06fF
C1698 s0 Gnd 36.69fF
C1699 b1out_1 Gnd 3.47fF
C1700 4bitadder_1/XOR_1/w_62_n20# Gnd 0.87fF
C1701 4bitadder_1/XOR_1/w_16_n1# Gnd 0.75fF
C1702 4bitadder_1/XOR_1/w_n34_n1# Gnd 0.75fF
C1703 4bitadder_1/XOR_1/w_62_37# Gnd 0.72fF
C1704 4bitadder_1/XOR_0/abar Gnd 0.12fF
C1705 4bitadder_1/XOR_0/bbar Gnd 0.06fF
C1706 b0out_1 Gnd 3.02fF
C1707 4bitadder_1/XOR_0/w_62_n20# Gnd 0.87fF
C1708 4bitadder_1/XOR_0/w_16_n1# Gnd 0.75fF
C1709 4bitadder_1/XOR_0/w_n34_n1# Gnd 0.75fF
C1710 4bitadder_1/XOR_0/w_62_37# Gnd 0.72fF
C1711 4bitadder_1/fulladder_3/XOR_1/abar Gnd 0.11fF
C1712 4bitadder_1/fulladder_3/XOR_1/bbar Gnd 0.06fF
C1713 s3_sub Gnd 1.05fF
C1714 4bitadder_1/fulladder_3/XOR_1/w_62_n20# Gnd 0.87fF
C1715 4bitadder_1/fulladder_3/XOR_1/w_16_n1# Gnd 0.75fF
C1716 4bitadder_1/fulladder_3/XOR_1/w_n34_n1# Gnd 0.75fF
C1717 4bitadder_1/fulladder_3/XOR_1/w_62_37# Gnd 0.72fF
C1718 4bitadder_1/fulladder_3/or_0/b Gnd 2.26fF
C1719 4bitadder_1/fulladder_3/and_1/a_n26_14# Gnd 0.05fF
C1720 a3out_1 Gnd 7.67fF
C1721 4bitadder_1/fulladder_3/and_1/w_26_9# Gnd 0.82fF
C1722 4bitadder_1/fulladder_3/and_1/w_n43_8# Gnd 0.82fF
C1723 4bitadder_1/fulladder_3/XOR_0/abar Gnd 0.11fF
C1724 4bitadder_1/fulladder_3/XOR_0/bbar Gnd 0.06fF
C1725 4bitadder_1/fulladder_3/XOR_0/w_62_n20# Gnd 0.87fF
C1726 4bitadder_1/fulladder_3/XOR_0/w_16_n1# Gnd 0.75fF
C1727 4bitadder_1/fulladder_3/XOR_0/w_n34_n1# Gnd 0.75fF
C1728 4bitadder_1/fulladder_3/XOR_0/w_62_37# Gnd 0.72fF
C1729 4bitadder_1/fulladder_3/or_0/a Gnd 1.96fF
C1730 4bitadder_1/fulladder_3/and_0/a_n26_14# Gnd 0.05fF
C1731 4bitadder_1/c3 Gnd 2.24fF
C1732 4bitadder_1/fulladder_3/axorb Gnd 3.25fF
C1733 4bitadder_1/fulladder_3/and_0/w_26_9# Gnd 0.82fF
C1734 4bitadder_1/fulladder_3/and_0/w_n43_8# Gnd 0.82fF
C1735 fc_sub Gnd 0.60fF
C1736 4bitadder_1/fulladder_3/or_0/a_n15_32# Gnd 0.17fF
C1737 4bitadder_1/fulladder_3/or_0/w_58_101# Gnd 1.55fF
C1738 4bitadder_1/fulladder_3/or_0/w_n48_101# Gnd 2.56fF
C1739 4bitadder_1/fulladder_2/XOR_1/abar Gnd 0.11fF
C1740 4bitadder_1/fulladder_2/XOR_1/bbar Gnd 0.06fF
C1741 s2_sub Gnd 0.72fF
C1742 4bitadder_1/fulladder_2/XOR_1/w_62_n20# Gnd 0.87fF
C1743 4bitadder_1/fulladder_2/XOR_1/w_16_n1# Gnd 0.75fF
C1744 4bitadder_1/fulladder_2/XOR_1/w_n34_n1# Gnd 0.75fF
C1745 4bitadder_1/fulladder_2/XOR_1/w_62_37# Gnd 0.72fF
C1746 4bitadder_1/fulladder_2/or_0/b Gnd 2.26fF
C1747 4bitadder_1/fulladder_2/and_1/a_n26_14# Gnd 0.05fF
C1748 4bitadder_1/XOR_2/out Gnd 2.12fF
C1749 4bitadder_1/fulladder_2/and_1/w_26_9# Gnd 0.82fF
C1750 4bitadder_1/fulladder_2/and_1/w_n43_8# Gnd 0.82fF
C1751 4bitadder_1/fulladder_2/XOR_0/abar Gnd 0.11fF
C1752 4bitadder_1/fulladder_2/XOR_0/bbar Gnd 0.06fF
C1753 4bitadder_1/fulladder_2/XOR_0/w_62_n20# Gnd 0.87fF
C1754 4bitadder_1/fulladder_2/XOR_0/w_16_n1# Gnd 0.75fF
C1755 4bitadder_1/fulladder_2/XOR_0/w_n34_n1# Gnd 0.75fF
C1756 4bitadder_1/fulladder_2/XOR_0/w_62_37# Gnd 0.72fF
C1757 4bitadder_1/fulladder_2/or_0/a Gnd 1.96fF
C1758 4bitadder_1/fulladder_2/and_0/a_n26_14# Gnd 0.05fF
C1759 4bitadder_1/fulladder_2/axorb Gnd 3.25fF
C1760 4bitadder_1/fulladder_2/and_0/w_26_9# Gnd 0.82fF
C1761 4bitadder_1/fulladder_2/and_0/w_n43_8# Gnd 0.82fF
C1762 4bitadder_1/fulladder_2/or_0/a_n15_32# Gnd 0.17fF
C1763 4bitadder_1/fulladder_2/or_0/w_58_101# Gnd 1.55fF
C1764 4bitadder_1/fulladder_2/or_0/w_n48_101# Gnd 2.56fF
C1765 4bitadder_1/fulladder_1/XOR_1/abar Gnd 0.11fF
C1766 4bitadder_1/fulladder_1/XOR_1/bbar Gnd 0.06fF
C1767 s1_sub Gnd 1.01fF
C1768 4bitadder_1/fulladder_1/XOR_1/w_62_n20# Gnd 0.87fF
C1769 4bitadder_1/fulladder_1/XOR_1/w_16_n1# Gnd 0.75fF
C1770 4bitadder_1/fulladder_1/XOR_1/w_n34_n1# Gnd 0.75fF
C1771 4bitadder_1/fulladder_1/XOR_1/w_62_37# Gnd 0.72fF
C1772 4bitadder_1/fulladder_1/or_0/b Gnd 2.26fF
C1773 4bitadder_1/fulladder_1/and_1/a_n26_14# Gnd 0.05fF
C1774 4bitadder_1/XOR_1/out Gnd 2.08fF
C1775 4bitadder_1/fulladder_1/and_1/w_26_9# Gnd 0.82fF
C1776 4bitadder_1/fulladder_1/and_1/w_n43_8# Gnd 0.82fF
C1777 4bitadder_1/fulladder_1/XOR_0/abar Gnd 0.11fF
C1778 4bitadder_1/fulladder_1/XOR_0/bbar Gnd 0.06fF
C1779 4bitadder_1/fulladder_1/XOR_0/w_62_n20# Gnd 0.87fF
C1780 4bitadder_1/fulladder_1/XOR_0/w_16_n1# Gnd 0.75fF
C1781 4bitadder_1/fulladder_1/XOR_0/w_n34_n1# Gnd 0.75fF
C1782 4bitadder_1/fulladder_1/XOR_0/w_62_37# Gnd 0.72fF
C1783 4bitadder_1/fulladder_1/or_0/a Gnd 1.96fF
C1784 4bitadder_1/fulladder_1/and_0/a_n26_14# Gnd 0.05fF
C1785 4bitadder_1/fulladder_1/axorb Gnd 3.25fF
C1786 4bitadder_1/fulladder_1/and_0/w_26_9# Gnd 0.82fF
C1787 4bitadder_1/fulladder_1/and_0/w_n43_8# Gnd 0.82fF
C1788 4bitadder_1/fulladder_1/or_0/a_n15_32# Gnd 0.17fF
C1789 4bitadder_1/fulladder_1/or_0/w_58_101# Gnd 1.55fF
C1790 4bitadder_1/fulladder_1/or_0/w_n48_101# Gnd 2.56fF
C1791 4bitadder_1/fulladder_0/XOR_1/abar Gnd 0.11fF
C1792 4bitadder_1/fulladder_0/XOR_1/bbar Gnd 0.06fF
C1793 s0_sub Gnd 0.46fF
C1794 4bitadder_1/fulladder_0/XOR_1/w_62_n20# Gnd 0.87fF
C1795 4bitadder_1/fulladder_0/XOR_1/w_16_n1# Gnd 0.75fF
C1796 4bitadder_1/fulladder_0/XOR_1/w_n34_n1# Gnd 0.75fF
C1797 4bitadder_1/fulladder_0/XOR_1/w_62_37# Gnd 0.72fF
C1798 4bitadder_1/fulladder_0/or_0/b Gnd 2.26fF
C1799 4bitadder_1/fulladder_0/and_1/a_n26_14# Gnd 0.05fF
C1800 a0_out1 Gnd 7.61fF
C1801 4bitadder_1/b0xorM Gnd 2.11fF
C1802 4bitadder_1/fulladder_0/and_1/w_26_9# Gnd 0.82fF
C1803 4bitadder_1/fulladder_0/and_1/w_n43_8# Gnd 0.82fF
C1804 4bitadder_1/fulladder_0/XOR_0/abar Gnd 0.11fF
C1805 4bitadder_1/fulladder_0/XOR_0/bbar Gnd 0.06fF
C1806 4bitadder_1/fulladder_0/XOR_0/w_62_n20# Gnd 0.87fF
C1807 4bitadder_1/fulladder_0/XOR_0/w_16_n1# Gnd 0.75fF
C1808 4bitadder_1/fulladder_0/XOR_0/w_n34_n1# Gnd 0.75fF
C1809 4bitadder_1/fulladder_0/XOR_0/w_62_37# Gnd 0.72fF
C1810 4bitadder_1/fulladder_0/or_0/a Gnd 1.96fF
C1811 4bitadder_1/fulladder_0/and_0/a_n26_14# Gnd 0.05fF
C1812 4bitadder_1/fulladder_0/axorb Gnd 3.25fF
C1813 4bitadder_1/fulladder_0/and_0/w_26_9# Gnd 0.82fF
C1814 4bitadder_1/fulladder_0/and_0/w_n43_8# Gnd 0.82fF
C1815 4bitadder_1/fulladder_0/or_0/a_n15_32# Gnd 0.17fF
C1816 4bitadder_1/fulladder_0/or_0/w_58_101# Gnd 1.55fF
C1817 4bitadder_1/fulladder_0/or_0/w_n48_101# Gnd 2.56fF
C1818 comparator_0/a2bar Gnd 5.34fF
C1819 comparator_0/3input_AND_1/w_69_n71# Gnd 1.13fF
C1820 comparator_0/3input_AND_1/w_32_n21# Gnd 1.13fF
C1821 comparator_0/3input_AND_1/w_n14_24# Gnd 1.13fF
C1822 gnd Gnd 99.11fF
C1823 comparator_0/t2 Gnd 3.00fF
C1824 comparator_0/3input_AND_1/not_0/in Gnd 1.59fF
C1825 comparator_0/3input_AND_1/not_0/w_n2_10# Gnd 0.90fF
C1826 comparator_0/b2bar Gnd 5.92fF
C1827 comparator_0/3input_AND_0/w_69_n71# Gnd 1.13fF
C1828 comparator_0/3input_AND_0/w_32_n21# Gnd 1.13fF
C1829 comparator_0/3input_AND_0/w_n14_24# Gnd 1.13fF
C1830 comparator_0/t6 Gnd 2.94fF
C1831 comparator_0/3input_AND_0/not_0/in Gnd 1.59fF
C1832 comparator_0/3input_AND_0/not_0/w_n2_10# Gnd 0.90fF
C1833 comparator_0/a2xnorb2 Gnd 18.99fF
C1834 comparator_0/4input_AND_2/w_68_n95# Gnd 1.13fF
C1835 comparator_0/4input_AND_2/w_29_n46# Gnd 1.13fF
C1836 comparator_0/4input_AND_2/w_n8_2# Gnd 1.13fF
C1837 comparator_0/4input_AND_2/w_n47_52# Gnd 1.13fF
C1838 comparator_0/t3 Gnd 4.44fF
C1839 comparator_0/4input_AND_2/not_0/in Gnd 2.38fF
C1840 comparator_0/4input_AND_2/not_0/w_n2_10# Gnd 0.90fF
C1841 comparator_0/and_1/a_n26_14# Gnd 0.05fF
C1842 comparator_0/a3bar Gnd 4.39fF
C1843 comparator_0/and_1/w_26_9# Gnd 0.82fF
C1844 comparator_0/and_1/w_n43_8# Gnd 0.82fF
C1845 comparator_0/4input_AND_1/w_68_n95# Gnd 1.13fF
C1846 comparator_0/4input_AND_1/w_29_n46# Gnd 1.13fF
C1847 comparator_0/4input_AND_1/w_n8_2# Gnd 1.13fF
C1848 comparator_0/4input_AND_1/w_n47_52# Gnd 1.13fF
C1849 comparator_0/t7 Gnd 4.39fF
C1850 comparator_0/4input_AND_1/not_0/in Gnd 2.38fF
C1851 comparator_0/4input_AND_1/not_0/w_n2_10# Gnd 0.90fF
C1852 comparator_0/4input_AND_0/w_68_n95# Gnd 1.13fF
C1853 comparator_0/4input_AND_0/w_29_n46# Gnd 1.13fF
C1854 comparator_0/4input_AND_0/w_n8_2# Gnd 1.13fF
C1855 comparator_0/4input_AND_0/w_n47_52# Gnd 1.13fF
C1856 equal Gnd 0.22fF
C1857 comparator_0/4input_AND_0/not_0/in Gnd 2.38fF
C1858 comparator_0/4input_AND_0/not_0/w_n2_10# Gnd 0.90fF
C1859 comparator_0/and_0/a_n26_14# Gnd 0.05fF
C1860 comparator_0/b3bar Gnd 0.68fF
C1861 comparator_0/and_0/w_26_9# Gnd 0.82fF
C1862 comparator_0/and_0/w_n43_8# Gnd 0.82fF
C1863 comparator_0/5input_AND_1/w_106_n113# Gnd 0.81fF
C1864 comparator_0/5input_AND_1/w_68_n82# Gnd 0.81fF
C1865 comparator_0/5input_AND_1/w_31_n55# Gnd 1.18fF
C1866 comparator_0/5input_AND_1/w_n4_n20# Gnd 0.89fF
C1867 comparator_0/5input_AND_1/w_n37_15# Gnd 0.89fF
C1868 comparator_0/t4 Gnd 2.77fF
C1869 comparator_0/5input_AND_1/not_0/in Gnd 2.73fF
C1870 comparator_0/5input_AND_1/not_0/w_n2_10# Gnd 0.90fF
C1871 comparator_0/5input_AND_0/w_106_n113# Gnd 0.81fF
C1872 comparator_0/5input_AND_0/w_68_n82# Gnd 0.81fF
C1873 comparator_0/5input_AND_0/w_31_n55# Gnd 1.18fF
C1874 comparator_0/5input_AND_0/w_n4_n20# Gnd 0.89fF
C1875 comparator_0/5input_AND_0/w_n37_15# Gnd 0.89fF
C1876 comparator_0/t8 Gnd 1.96fF
C1877 comparator_0/5input_AND_0/not_0/in Gnd 2.73fF
C1878 comparator_0/5input_AND_0/not_0/w_n2_10# Gnd 0.90fF
C1879 comparator_0/not_7/w_n2_10# Gnd 0.90fF
C1880 comparator_0/not_6/w_n2_10# Gnd 0.90fF
C1881 comparator_0/a1bar Gnd 5.03fF
C1882 comparator_0/not_5/w_n2_10# Gnd 0.90fF
C1883 comparator_0/xnor_3/XOR_0/abar Gnd 0.11fF
C1884 comparator_0/xnor_3/XOR_0/bbar Gnd 0.06fF
C1885 comparator_0/xnor_3/not_0/in Gnd 0.39fF
C1886 boout_2 Gnd 8.80fF
C1887 a0out_2 Gnd 32.03fF
C1888 comparator_0/xnor_3/XOR_0/w_62_n20# Gnd 0.87fF
C1889 comparator_0/xnor_3/XOR_0/w_16_n1# Gnd 0.75fF
C1890 comparator_0/xnor_3/XOR_0/w_n34_n1# Gnd 0.75fF
C1891 comparator_0/xnor_3/XOR_0/w_62_37# Gnd 0.72fF
C1892 comparator_0/a0xnorb0 Gnd 2.96fF
C1893 comparator_0/xnor_3/not_0/w_n2_10# Gnd 0.90fF
C1894 comparator_0/xnor_2/XOR_0/abar Gnd 0.11fF
C1895 comparator_0/xnor_2/XOR_0/bbar Gnd 0.06fF
C1896 comparator_0/xnor_2/not_0/in Gnd 0.39fF
C1897 b1out_2 Gnd 55.09fF
C1898 a1out_2 Gnd 41.81fF
C1899 comparator_0/xnor_2/XOR_0/w_62_n20# Gnd 0.87fF
C1900 comparator_0/xnor_2/XOR_0/w_16_n1# Gnd 0.75fF
C1901 comparator_0/xnor_2/XOR_0/w_n34_n1# Gnd 0.75fF
C1902 comparator_0/xnor_2/XOR_0/w_62_37# Gnd 0.72fF
C1903 comparator_0/xnor_2/not_0/w_n2_10# Gnd 0.90fF
C1904 comparator_0/4input_OR_1/w_n58_n43# Gnd 2.55fF
C1905 bga Gnd 0.14fF
C1906 comparator_0/4input_OR_1/y Gnd 1.46fF
C1907 comparator_0/4input_OR_1/NOT_0/w_n2_10# Gnd 0.90fF
C1908 comparator_0/a0bar Gnd 6.16fF
C1909 comparator_0/not_4/w_n2_10# Gnd 0.90fF
C1910 comparator_0/xnor_1/XOR_0/abar Gnd 0.11fF
C1911 comparator_0/xnor_1/XOR_0/bbar Gnd 0.06fF
C1912 comparator_0/xnor_1/not_0/in Gnd 0.39fF
C1913 b2out_2 Gnd 46.65fF
C1914 a2out_2 Gnd 27.86fF
C1915 comparator_0/xnor_1/XOR_0/w_62_n20# Gnd 0.87fF
C1916 comparator_0/xnor_1/XOR_0/w_16_n1# Gnd 0.75fF
C1917 comparator_0/xnor_1/XOR_0/w_n34_n1# Gnd 0.75fF
C1918 comparator_0/xnor_1/XOR_0/w_62_37# Gnd 0.72fF
C1919 comparator_0/xnor_1/not_0/w_n2_10# Gnd 0.90fF
C1920 comparator_0/not_3/w_n2_10# Gnd 0.90fF
C1921 comparator_0/xnor_0/XOR_0/abar Gnd 0.11fF
C1922 comparator_0/xnor_0/XOR_0/bbar Gnd 0.06fF
C1923 comparator_0/xnor_0/not_0/in Gnd 0.39fF
C1924 comparator_0/b3 Gnd 44.13fF
C1925 a3out_2 Gnd 20.89fF
C1926 comparator_0/xnor_0/XOR_0/w_62_n20# Gnd 0.87fF
C1927 comparator_0/xnor_0/XOR_0/w_16_n1# Gnd 0.75fF
C1928 comparator_0/xnor_0/XOR_0/w_n34_n1# Gnd 0.75fF
C1929 comparator_0/xnor_0/XOR_0/w_62_37# Gnd 0.72fF
C1930 comparator_0/xnor_0/not_0/w_n2_10# Gnd 0.90fF
C1931 comparator_0/not_2/w_n2_10# Gnd 0.90fF
C1932 comparator_0/4input_OR_0/w_n58_n43# Gnd 2.55fF
C1933 agb Gnd 0.14fF
C1934 comparator_0/4input_OR_0/y Gnd 1.46fF
C1935 vdd Gnd 121.02fF
C1936 comparator_0/4input_OR_0/NOT_0/w_n2_10# Gnd 0.90fF
C1937 comparator_0/b1bar Gnd 4.66fF
C1938 comparator_0/not_1/w_n2_10# Gnd 0.90fF
C1939 comparator_0/b0bar Gnd 6.97fF
C1940 comparator_0/not_0/w_n2_10# Gnd 0.90fF
C1941 4bitadder_0/XOR_3/abar Gnd 0.11fF
C1942 4bitadder_0/XOR_3/bbar Gnd 0.06fF
C1943 4bitadder_0/XOR_3/w_62_n20# Gnd 0.87fF
C1944 4bitadder_0/XOR_3/w_16_n1# Gnd 0.75fF
C1945 4bitadder_0/XOR_3/w_n34_n1# Gnd 0.75fF
C1946 4bitadder_0/XOR_3/w_62_37# Gnd 0.72fF
C1947 4bitadder_0/XOR_2/abar Gnd 0.11fF
C1948 4bitadder_0/XOR_2/bbar Gnd 0.06fF
C1949 4bitadder_0/XOR_2/w_62_n20# Gnd 0.87fF
C1950 4bitadder_0/XOR_2/w_16_n1# Gnd 0.75fF
C1951 4bitadder_0/XOR_2/w_n34_n1# Gnd 0.75fF
C1952 4bitadder_0/XOR_2/w_62_37# Gnd 0.72fF
C1953 4bitadder_0/XOR_1/abar Gnd 0.11fF
C1954 4bitadder_0/XOR_1/bbar Gnd 0.06fF
C1955 4bitadder_0/XOR_1/w_62_n20# Gnd 0.87fF
C1956 4bitadder_0/XOR_1/w_16_n1# Gnd 0.75fF
C1957 4bitadder_0/XOR_1/w_n34_n1# Gnd 0.75fF
C1958 4bitadder_0/XOR_1/w_62_37# Gnd 0.72fF
C1959 4bitadder_0/XOR_0/abar Gnd 0.12fF
C1960 4bitadder_0/XOR_0/bbar Gnd 0.06fF
C1961 4bitadder_0/XOR_0/w_62_n20# Gnd 0.87fF
C1962 4bitadder_0/XOR_0/w_16_n1# Gnd 0.75fF
C1963 4bitadder_0/XOR_0/w_n34_n1# Gnd 0.75fF
C1964 4bitadder_0/XOR_0/w_62_37# Gnd 0.72fF
C1965 4bitadder_0/fulladder_3/XOR_1/abar Gnd 0.11fF
C1966 4bitadder_0/fulladder_3/XOR_1/bbar Gnd 0.06fF
C1967 s3_add Gnd 0.74fF
C1968 4bitadder_0/fulladder_3/XOR_1/w_62_n20# Gnd 0.87fF
C1969 4bitadder_0/fulladder_3/XOR_1/w_16_n1# Gnd 0.75fF
C1970 4bitadder_0/fulladder_3/XOR_1/w_n34_n1# Gnd 0.75fF
C1971 4bitadder_0/fulladder_3/XOR_1/w_62_37# Gnd 0.72fF
C1972 4bitadder_0/fulladder_3/or_0/b Gnd 2.26fF
C1973 4bitadder_0/fulladder_3/and_1/a_n26_14# Gnd 0.05fF
C1974 a3out_0 Gnd 7.66fF
C1975 4bitadder_0/fulladder_3/and_1/w_26_9# Gnd 0.82fF
C1976 4bitadder_0/fulladder_3/and_1/w_n43_8# Gnd 0.82fF
C1977 4bitadder_0/fulladder_3/XOR_0/abar Gnd 0.11fF
C1978 4bitadder_0/fulladder_3/XOR_0/bbar Gnd 0.06fF
C1979 4bitadder_0/fulladder_3/XOR_0/w_62_n20# Gnd 0.87fF
C1980 4bitadder_0/fulladder_3/XOR_0/w_16_n1# Gnd 0.75fF
C1981 4bitadder_0/fulladder_3/XOR_0/w_n34_n1# Gnd 0.75fF
C1982 4bitadder_0/fulladder_3/XOR_0/w_62_37# Gnd 0.72fF
C1983 4bitadder_0/fulladder_3/or_0/a Gnd 1.96fF
C1984 4bitadder_0/fulladder_3/and_0/a_n26_14# Gnd 0.05fF
C1985 4bitadder_0/c3 Gnd 2.24fF
C1986 4bitadder_0/fulladder_3/axorb Gnd 3.25fF
C1987 4bitadder_0/fulladder_3/and_0/w_26_9# Gnd 0.82fF
C1988 4bitadder_0/fulladder_3/and_0/w_n43_8# Gnd 0.82fF
C1989 fc_add Gnd 0.54fF
C1990 4bitadder_0/fulladder_3/or_0/a_n15_32# Gnd 0.17fF
C1991 4bitadder_0/fulladder_3/or_0/w_58_101# Gnd 1.55fF
C1992 4bitadder_0/fulladder_3/or_0/w_n48_101# Gnd 2.56fF
C1993 4bitadder_0/fulladder_2/XOR_1/abar Gnd 0.11fF
C1994 4bitadder_0/fulladder_2/XOR_1/bbar Gnd 0.06fF
C1995 s2_add Gnd 0.65fF
C1996 4bitadder_0/fulladder_2/XOR_1/w_62_n20# Gnd 0.87fF
C1997 4bitadder_0/fulladder_2/XOR_1/w_16_n1# Gnd 0.75fF
C1998 4bitadder_0/fulladder_2/XOR_1/w_n34_n1# Gnd 0.75fF
C1999 4bitadder_0/fulladder_2/XOR_1/w_62_37# Gnd 0.72fF
C2000 4bitadder_0/fulladder_2/or_0/b Gnd 2.26fF
C2001 4bitadder_0/fulladder_2/and_1/a_n26_14# Gnd 0.05fF
C2002 a2out_0 Gnd 7.81fF
C2003 4bitadder_0/XOR_2/out Gnd 2.12fF
C2004 4bitadder_0/fulladder_2/and_1/w_26_9# Gnd 0.82fF
C2005 4bitadder_0/fulladder_2/and_1/w_n43_8# Gnd 0.82fF
C2006 4bitadder_0/fulladder_2/XOR_0/abar Gnd 0.11fF
C2007 4bitadder_0/fulladder_2/XOR_0/bbar Gnd 0.06fF
C2008 4bitadder_0/fulladder_2/XOR_0/w_62_n20# Gnd 0.87fF
C2009 4bitadder_0/fulladder_2/XOR_0/w_16_n1# Gnd 0.75fF
C2010 4bitadder_0/fulladder_2/XOR_0/w_n34_n1# Gnd 0.75fF
C2011 4bitadder_0/fulladder_2/XOR_0/w_62_37# Gnd 0.72fF
C2012 4bitadder_0/fulladder_2/or_0/a Gnd 1.96fF
C2013 4bitadder_0/fulladder_2/and_0/a_n26_14# Gnd 0.05fF
C2014 4bitadder_0/fulladder_2/axorb Gnd 3.25fF
C2015 4bitadder_0/fulladder_2/and_0/w_26_9# Gnd 0.82fF
C2016 4bitadder_0/fulladder_2/and_0/w_n43_8# Gnd 0.82fF
C2017 4bitadder_0/fulladder_2/or_0/a_n15_32# Gnd 0.17fF
C2018 4bitadder_0/fulladder_2/or_0/w_58_101# Gnd 1.55fF
C2019 4bitadder_0/fulladder_2/or_0/w_n48_101# Gnd 2.56fF
C2020 4bitadder_0/fulladder_1/XOR_1/abar Gnd 0.11fF
C2021 4bitadder_0/fulladder_1/XOR_1/bbar Gnd 0.06fF
C2022 s1_add Gnd 1.15fF
C2023 4bitadder_0/fulladder_1/XOR_1/w_62_n20# Gnd 0.87fF
C2024 4bitadder_0/fulladder_1/XOR_1/w_16_n1# Gnd 0.75fF
C2025 4bitadder_0/fulladder_1/XOR_1/w_n34_n1# Gnd 0.75fF
C2026 4bitadder_0/fulladder_1/XOR_1/w_62_37# Gnd 0.72fF
C2027 4bitadder_0/fulladder_1/or_0/b Gnd 2.26fF
C2028 4bitadder_0/fulladder_1/and_1/a_n26_14# Gnd 0.05fF
C2029 a1out_0 Gnd 7.72fF
C2030 4bitadder_0/XOR_1/out Gnd 2.08fF
C2031 4bitadder_0/fulladder_1/and_1/w_26_9# Gnd 0.82fF
C2032 4bitadder_0/fulladder_1/and_1/w_n43_8# Gnd 0.82fF
C2033 4bitadder_0/fulladder_1/XOR_0/abar Gnd 0.11fF
C2034 4bitadder_0/fulladder_1/XOR_0/bbar Gnd 0.06fF
C2035 4bitadder_0/fulladder_1/XOR_0/w_62_n20# Gnd 0.87fF
C2036 4bitadder_0/fulladder_1/XOR_0/w_16_n1# Gnd 0.75fF
C2037 4bitadder_0/fulladder_1/XOR_0/w_n34_n1# Gnd 0.75fF
C2038 4bitadder_0/fulladder_1/XOR_0/w_62_37# Gnd 0.72fF
C2039 4bitadder_0/fulladder_1/or_0/a Gnd 1.96fF
C2040 4bitadder_0/fulladder_1/and_0/a_n26_14# Gnd 0.05fF
C2041 4bitadder_0/fulladder_1/axorb Gnd 3.25fF
C2042 4bitadder_0/fulladder_1/and_0/w_26_9# Gnd 0.82fF
C2043 4bitadder_0/fulladder_1/and_0/w_n43_8# Gnd 0.82fF
C2044 4bitadder_0/fulladder_1/or_0/a_n15_32# Gnd 0.17fF
C2045 4bitadder_0/fulladder_1/or_0/w_58_101# Gnd 1.55fF
C2046 4bitadder_0/fulladder_1/or_0/w_n48_101# Gnd 2.56fF
C2047 4bitadder_0/fulladder_0/XOR_1/abar Gnd 0.11fF
C2048 4bitadder_0/fulladder_0/XOR_1/bbar Gnd 0.06fF
C2049 s0_add Gnd 0.87fF
C2050 4bitadder_0/fulladder_0/XOR_1/w_62_n20# Gnd 0.87fF
C2051 4bitadder_0/fulladder_0/XOR_1/w_16_n1# Gnd 0.75fF
C2052 4bitadder_0/fulladder_0/XOR_1/w_n34_n1# Gnd 0.75fF
C2053 4bitadder_0/fulladder_0/XOR_1/w_62_37# Gnd 0.72fF
C2054 4bitadder_0/fulladder_0/or_0/b Gnd 2.26fF
C2055 4bitadder_0/fulladder_0/and_1/a_n26_14# Gnd 0.05fF
C2056 a0out_0 Gnd 7.55fF
C2057 4bitadder_0/b0xorM Gnd 2.11fF
C2058 4bitadder_0/fulladder_0/and_1/w_26_9# Gnd 0.82fF
C2059 4bitadder_0/fulladder_0/and_1/w_n43_8# Gnd 0.82fF
C2060 4bitadder_0/fulladder_0/XOR_0/abar Gnd 0.11fF
C2061 4bitadder_0/fulladder_0/XOR_0/bbar Gnd 0.06fF
C2062 4bitadder_0/fulladder_0/XOR_0/w_62_n20# Gnd 0.87fF
C2063 4bitadder_0/fulladder_0/XOR_0/w_16_n1# Gnd 0.75fF
C2064 4bitadder_0/fulladder_0/XOR_0/w_n34_n1# Gnd 0.75fF
C2065 4bitadder_0/fulladder_0/XOR_0/w_62_37# Gnd 0.72fF
C2066 4bitadder_0/fulladder_0/or_0/a Gnd 1.96fF
C2067 4bitadder_0/fulladder_0/and_0/a_n26_14# Gnd 0.05fF
C2068 4bitadder_0/fulladder_0/axorb Gnd 3.25fF
C2069 4bitadder_0/fulladder_0/and_0/w_26_9# Gnd 0.82fF
C2070 4bitadder_0/fulladder_0/and_0/w_n43_8# Gnd 0.82fF
C2071 4bitadder_0/fulladder_0/or_0/a_n15_32# Gnd 0.17fF
C2072 4bitadder_0/fulladder_0/or_0/w_58_101# Gnd 1.55fF
C2073 4bitadder_0/fulladder_0/or_0/w_n48_101# Gnd 2.56fF
C2074 out3 Gnd 0.20fF
C2075 AND_Block_0/and_3/a_n26_14# Gnd 0.05fF
C2076 b3out_3 Gnd 0.73fF
C2077 a3out_3 Gnd 0.75fF
C2078 AND_Block_0/and_3/w_26_9# Gnd 0.82fF
C2079 AND_Block_0/and_3/w_n43_8# Gnd 0.82fF
C2080 out2 Gnd 0.20fF
C2081 AND_Block_0/and_2/a_n26_14# Gnd 0.05fF
C2082 b2out_3 Gnd 0.74fF
C2083 a2out_3 Gnd 0.77fF
C2084 AND_Block_0/and_2/w_26_9# Gnd 0.82fF
C2085 AND_Block_0/and_2/w_n43_8# Gnd 0.82fF
C2086 out1 Gnd 0.21fF
C2087 AND_Block_0/and_1/a_n26_14# Gnd 0.05fF
C2088 b1out_3 Gnd 0.75fF
C2089 a1out_3 Gnd 0.79fF
C2090 AND_Block_0/and_1/w_26_9# Gnd 0.82fF
C2091 AND_Block_0/and_1/w_n43_8# Gnd 0.82fF
C2092 out0 Gnd 0.20fF
C2093 AND_Block_0/and_0/a_n26_14# Gnd 0.05fF
C2094 b0out_3 Gnd 0.72fF
C2095 AND_Block_0/and_0/w_26_9# Gnd 0.82fF
C2096 AND_Block_0/and_0/w_n43_8# Gnd 0.82fF
C2097 enable_2/and_4/a_n26_14# Gnd 0.05fF
C2098 enable_2/and_4/w_26_9# Gnd 0.82fF
C2099 enable_2/and_4/w_n43_8# Gnd 0.82fF
C2100 enable_2/and_3/a_n26_14# Gnd 0.05fF
C2101 enable_2/and_3/w_26_9# Gnd 0.82fF
C2102 enable_2/and_3/w_n43_8# Gnd 0.82fF
C2103 enable_2/and_2/a_n26_14# Gnd 0.05fF
C2104 enable_2/a2 Gnd 0.55fF
C2105 enable_2/and_2/w_26_9# Gnd 0.82fF
C2106 enable_2/and_2/w_n43_8# Gnd 0.82fF
C2107 enable_2/and_1/a_n26_14# Gnd 0.05fF
C2108 enable_2/and_1/w_26_9# Gnd 0.82fF
C2109 enable_2/and_1/w_n43_8# Gnd 0.82fF
C2110 enable_2/and_0/a_n26_14# Gnd 0.05fF
C2111 enable_2/a0 Gnd 0.55fF
C2112 enable_2/and_0/w_26_9# Gnd 0.82fF
C2113 enable_2/and_0/w_n43_8# Gnd 0.82fF
C2114 enable_2/and_6/a_n26_14# Gnd 0.05fF
C2115 enable_2/and_6/w_26_9# Gnd 0.82fF
C2116 enable_2/and_6/w_n43_8# Gnd 0.82fF
C2117 b3out_2 Gnd 0.40fF
C2118 enable_2/and_7/a_n26_14# Gnd 0.05fF
C2119 enable_2/en Gnd 2.76fF
C2120 enable_2/and_7/w_26_9# Gnd 0.82fF
C2121 enable_2/and_7/w_n43_8# Gnd 0.82fF
C2122 enable_2/and_5/a_n26_14# Gnd 0.05fF
C2123 enable_2/and_5/w_26_9# Gnd 0.82fF
C2124 enable_2/and_5/w_n43_8# Gnd 0.82fF
C2125 enable_3/and_4/a_n26_14# Gnd 0.05fF
C2126 b0 Gnd 1.59fF
C2127 enable_3/and_4/w_26_9# Gnd 0.82fF
C2128 enable_3/and_4/w_n43_8# Gnd 0.82fF
C2129 enable_3/and_3/a_n26_14# Gnd 0.05fF
C2130 a3 Gnd 1.58fF
C2131 enable_3/and_3/w_26_9# Gnd 0.82fF
C2132 enable_3/and_3/w_n43_8# Gnd 0.82fF
C2133 enable_3/and_2/a_n26_14# Gnd 0.05fF
C2134 a2 Gnd 1.18fF
C2135 enable_3/and_2/w_26_9# Gnd 0.82fF
C2136 enable_3/and_2/w_n43_8# Gnd 0.82fF
C2137 enable_3/and_1/a_n26_14# Gnd 0.05fF
C2138 enable_3/and_1/w_26_9# Gnd 0.82fF
C2139 enable_3/and_1/w_n43_8# Gnd 0.82fF
C2140 enable_3/and_0/a_n26_14# Gnd 0.05fF
C2141 a0 Gnd 1.17fF
C2142 enable_3/and_0/w_26_9# Gnd 0.82fF
C2143 enable_3/and_0/w_n43_8# Gnd 0.82fF
C2144 enable_3/and_6/a_n26_14# Gnd 0.05fF
C2145 b2 Gnd 1.57fF
C2146 enable_3/and_6/w_26_9# Gnd 0.82fF
C2147 enable_3/and_6/w_n43_8# Gnd 0.82fF
C2148 enable_3/and_7/a_n26_14# Gnd 0.05fF
C2149 b3 Gnd 1.60fF
C2150 enable_3/en Gnd 7.29fF
C2151 enable_3/and_7/w_26_9# Gnd 0.82fF
C2152 enable_3/and_7/w_n43_8# Gnd 0.82fF
C2153 enable_3/and_5/a_n26_14# Gnd 0.05fF
C2154 b1 Gnd 1.17fF
C2155 enable_3/and_5/w_26_9# Gnd 0.82fF
C2156 enable_3/and_5/w_n43_8# Gnd 0.82fF
C2157 enable_1/and_4/a_n26_14# Gnd 0.05fF
C2158 enable_1/and_4/w_26_9# Gnd 0.82fF
C2159 enable_1/and_4/w_n43_8# Gnd 0.82fF
C2160 enable_1/and_3/a_n26_14# Gnd 0.05fF
C2161 enable_1/and_3/w_26_9# Gnd 0.82fF
C2162 enable_1/and_3/w_n43_8# Gnd 0.82fF
C2163 enable_1/and_2/a_n26_14# Gnd 0.05fF
C2164 enable_1/and_2/w_26_9# Gnd 0.82fF
C2165 enable_1/and_2/w_n43_8# Gnd 0.82fF
C2166 enable_1/and_1/a_n26_14# Gnd 0.05fF
C2167 enable_1/and_1/w_26_9# Gnd 0.82fF
C2168 enable_1/and_1/w_n43_8# Gnd 0.82fF
C2169 enable_1/and_0/a_n26_14# Gnd 0.05fF
C2170 enable_1/and_0/w_26_9# Gnd 0.82fF
C2171 enable_1/and_0/w_n43_8# Gnd 0.82fF
C2172 enable_1/and_6/a_n26_14# Gnd 0.05fF
C2173 enable_1/and_6/w_26_9# Gnd 0.82fF
C2174 enable_1/and_6/w_n43_8# Gnd 0.82fF
C2175 enable_1/and_7/a_n26_14# Gnd 0.05fF
C2176 enable_1/en Gnd 2.89fF
C2177 enable_1/and_7/w_26_9# Gnd 0.82fF
C2178 enable_1/and_7/w_n43_8# Gnd 0.82fF
C2179 enable_1/and_5/a_n26_14# Gnd 0.05fF
C2180 enable_1/and_5/w_26_9# Gnd 0.82fF
C2181 enable_1/and_5/w_n43_8# Gnd 0.82fF
C2182 b0out_0 Gnd 3.00fF
C2183 enable_0/and_4/a_n26_14# Gnd 0.05fF
C2184 enable_0/and_4/w_26_9# Gnd 0.82fF
C2185 enable_0/and_4/w_n43_8# Gnd 0.82fF
C2186 enable_0/and_3/a_n26_14# Gnd 0.05fF
C2187 enable_0/and_3/w_26_9# Gnd 0.82fF
C2188 enable_0/and_3/w_n43_8# Gnd 0.82fF
C2189 enable_0/and_2/a_n26_14# Gnd 0.05fF
C2190 enable_0/and_2/w_26_9# Gnd 0.82fF
C2191 enable_0/and_2/w_n43_8# Gnd 0.82fF
C2192 enable_0/and_1/a_n26_14# Gnd 0.05fF
C2193 enable_0/and_1/w_26_9# Gnd 0.82fF
C2194 enable_0/and_1/w_n43_8# Gnd 0.82fF
C2195 enable_0/and_0/a_n26_14# Gnd 0.05fF
C2196 enable_0/and_0/w_26_9# Gnd 0.82fF
C2197 enable_0/and_0/w_n43_8# Gnd 0.82fF
C2198 enable_0/and_6/a_n26_14# Gnd 0.05fF
C2199 enable_0/and_6/w_26_9# Gnd 0.82fF
C2200 enable_0/and_6/w_n43_8# Gnd 0.82fF
C2201 enable_0/and_7/a_n26_14# Gnd 0.05fF
C2202 enable_0/en Gnd 3.37fF
C2203 enable_0/and_7/w_26_9# Gnd 0.82fF
C2204 enable_0/and_7/w_n43_8# Gnd 0.82fF
C2205 b1out_0 Gnd 2.82fF
C2206 enable_0/and_5/a_n26_14# Gnd 0.05fF
C2207 enable_0/and_5/w_26_9# Gnd 0.82fF
C2208 enable_0/and_5/w_n43_8# Gnd 0.82fF

.tran 0.1n 500n

.measure tran trise 
+ TRIG v(b3) VAL = 'SUPPLY/2' RISE =1
+ TARG v(s2_add) VAL = 'SUPPLY/2' RISE =1 

.measure tran tfall 
+ TRIG v(b3) VAL = 'SUPPLY/2' FALL =1 
+ TARG v(s2_add) VAL = 'SUPPLY/2' FALL=1

.measure tran tpd param = '(trise + tfall)/2' goal = 0
        
.control
run
quit
* plot v(a0) v(a1)+2 v(a2)+4 v(a3)+6
* plot v(b0) v(b1)+2 v(b2)+4 v(b3)+6
* * plot v(a0out_3) v(a1out_3)+2 v(a2out_3)+4 v(a3out_3)+6
* * plot v(b0out_3) v(b1out_3)+2 v(b2out_3)+4 v(b3out_3)+6
* * plot v(s0_add) v(s1_add)+2 v(s2_add)+4 v(s3_add)+6 v(fc_add)+8
* * plot v(s0_sub) v(s1_sub)+2 v(s2_sub)+4 v(s3_sub)+6 v(fc_sub)+8
* plot v(out0) v(out1)+2 v(out2)+4 v(out3)+6

.endc

.end

