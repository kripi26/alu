* SPICE3 file created from xnor.ext - technology: scmos
.include TSMC_180nm.txt
.param SUPPLY = 1.8
.param LAMBDA = 0.09u
.param width_P = 8*LAMBDA
.param width_N = 4*LAMBDA
.global gnd vdd
.option scale=0.09u

Vdd vdd gnd 1.8
va a gnd pulse 0 1.8 0ns 100ps 100ps 60ns 100ns
vb b gnd pulse 0 1.8 0ns 100ps 100ps 20ns 60ns
.option scale=0.09u

M1000 y not_0/in vdd not_0/vdd CMOSP w=8 l=4
+  ad=101 pd=42 as=201 ps=102
M1001 y not_0/in gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=91 ps=40
M1002 not_0/in b XOR_0/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1003 XOR_0/bbar b XOR_0/gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=836 ps=164
M1004 not_0/in XOR_0/bbar XOR_0/abar XOR_0/vdd CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1005 vdd b XOR_0/bbar XOR_0/vdd CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1006 not_0/in b a XOR_0/vdd CMOSP w=8 l=6
+  ad=0 pd=0 as=72 ps=34
M1007 XOR_0/abar a XOR_0/gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1008 vdd a XOR_0/abar XOR_0/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1009 not_0/in XOR_0/bbar a Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=165 ps=52
C0 XOR_0/vdd XOR_0/bbar 0.03fF
C1 XOR_0/w_n34_n1# XOR_0/abar 0.03fF
C2 not_0/vdd not_0/in 0.09fF
C3 a XOR_0/w_n34_n1# 0.11fF
C4 vdd a 0.10fF
C5 XOR_0/abar b 0.30fF
C6 b XOR_0/gnd 0.33fF
C7 b not_0/in 0.13fF
C8 XOR_0/vdd not_0/in 0.02fF
C9 a XOR_0/vdd 0.02fF
C10 vdd not_0/vdd 0.18fF
C11 XOR_0/vdd XOR_0/bbar 0.13fF
C12 vdd XOR_0/w_n34_n1# 0.02fF
C13 not_0/vdd y 0.03fF
C14 vdd y 0.04fF
C15 vdd XOR_0/vdd 0.02fF
C16 XOR_0/vdd b 0.13fF
C17 XOR_0/abar gnd 0.07fF
C18 XOR_0/vdd XOR_0/abar 0.02fF
C19 a XOR_0/abar 0.13fF
C20 XOR_0/bbar b 0.02fF
C21 XOR_0/vdd b 0.11fF
C22 gnd XOR_0/gnd 0.07fF
C23 gnd not_0/in 0.03fF
C24 XOR_0/vdd not_0/in 0.04fF
C25 XOR_0/gnd Gnd 0.25fF
C26 XOR_0/abar Gnd 0.11fF
C27 XOR_0/bbar Gnd 0.06fF
C28 not_0/in Gnd 0.39fF
C29 b Gnd 1.52fF
C30 vdd Gnd 0.46fF
C31 a Gnd 2.79fF
C32 XOR_0/vdd Gnd 0.87fF
C33 XOR_0/vdd Gnd 0.75fF
C34 XOR_0/w_n34_n1# Gnd 0.75fF
C35 XOR_0/vdd Gnd 0.72fF
C36 gnd Gnd 0.62fF
C37 y Gnd 0.06fF
C38 not_0/vdd Gnd 0.90fF

.tran 0.1n 500n

* .measure tran trise
* + TRIG v(a) VAL = 0.9 RISE = 1
* + TARG v(out) VAL = 0.9 FALL = 1

* .measure tran tfall
* + TRIG v(a) VAL = 0.9 FALL = 1
* + TARG v(out) VAL = 0.9 RISE = 1

* .measure tran tpd param = '(trise + tfall)/2' goal = 0

.control
run
plot  v(a) v(b)+2 v(y)+4
.endc

.end


