* SPICE3 file created from alu.ext - technology: scmos
* SPICE3 file created from alu.ext - technology: scmos
.include TSMC_180nm.txt
.param SUPPLY = 1.8
.param LAMBDA = 0.09u
.param width_P = 8*LAMBDA
.param width_N = 4*LAMBDA
.global gnd vdd

Vdd vdd gnd 1.8
vs0 s0 gnd DC 0
vs1 s1 gnd DC 1.8
va0 a0 gnd pulse 0 1.8 0ns 100ps 100ps 20ns 40ns
va1 a1 gnd pulse 0 1.8 0ns 100ps 100ps 40ns 60ns
va2 a2 gnd pulse 0 1.8 0ns 100ps 100ps 60ns 80ns
va3 a3 gnd pulse 0 1.8 0ns 100ps 100ps 80ns 100ns
vb0 b0 gnd pulse 0 1.8 0ns 100ps 100ps 40ns 60ns
vb1 b1 gnd pulse 0 1.8 0ns 100ps 100ps 20ns 40ns
vb2 b2 gnd pulse 0 1.8 0ns 100ps 100ps 60ns 80ns
vb3 b3 gnd pulse 0 1.8 0ns 100ps 100ps 80ns 100ns

.option scale=0.09u

M1000 b1out_0 enable_0/and_5/a_n26_14# vdd enable_0/and_5/w_26_9# CMOSP w=7 l=4
+  ad=184 pd=80 as=24003 ps=10478
M1001 vdd b1 enable_0/and_5/a_n26_14# enable_0/and_5/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1002 b1out_0 enable_0/and_5/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=309 pd=102 as=48401 ps=12710
M1003 enable_0/and_5/a_n26_14# enable_0/en vdd enable_0/and_5/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1004 enable_0/and_5/a_n26_n23# enable_0/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1005 enable_0/and_5/a_n26_14# b1 enable_0/and_5/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1006 b3out_0 enable_0/and_7/a_n26_14# vdd enable_0/and_7/w_26_9# CMOSP w=7 l=4
+  ad=184 pd=80 as=0 ps=0
M1007 vdd b3 enable_0/and_7/a_n26_14# enable_0/and_7/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1008 b3out_0 enable_0/and_7/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=309 pd=102 as=0 ps=0
M1009 enable_0/and_7/a_n26_14# enable_0/en vdd enable_0/and_7/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1010 enable_0/and_7/a_n26_n23# enable_0/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1011 enable_0/and_7/a_n26_14# b3 enable_0/and_7/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1012 b2out_0 enable_0/and_6/a_n26_14# vdd enable_0/and_6/w_26_9# CMOSP w=7 l=4
+  ad=184 pd=80 as=0 ps=0
M1013 vdd b2 enable_0/and_6/a_n26_14# enable_0/and_6/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1014 b2out_0 enable_0/and_6/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=309 pd=102 as=0 ps=0
M1015 enable_0/and_6/a_n26_14# enable_0/en vdd enable_0/and_6/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1016 enable_0/and_6/a_n26_n23# enable_0/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1017 enable_0/and_6/a_n26_14# b2 enable_0/and_6/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1018 a0out_0 enable_0/and_0/a_n26_14# vdd enable_0/and_0/w_26_9# CMOSP w=7 l=4
+  ad=184 pd=80 as=0 ps=0
M1019 vdd a0 enable_0/and_0/a_n26_14# enable_0/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1020 a0out_0 enable_0/and_0/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=309 pd=102 as=0 ps=0
M1021 enable_0/and_0/a_n26_14# enable_0/en vdd enable_0/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1022 enable_0/and_0/a_n26_n23# enable_0/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1023 enable_0/and_0/a_n26_14# a0 enable_0/and_0/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1024 a1out_0 enable_0/and_1/a_n26_14# vdd enable_0/and_1/w_26_9# CMOSP w=7 l=4
+  ad=184 pd=80 as=0 ps=0
M1025 vdd a1 enable_0/and_1/a_n26_14# enable_0/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1026 a1out_0 enable_0/and_1/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=309 pd=102 as=0 ps=0
M1027 enable_0/and_1/a_n26_14# enable_0/en vdd enable_0/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1028 enable_0/and_1/a_n26_n23# enable_0/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1029 enable_0/and_1/a_n26_14# a1 enable_0/and_1/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1030 a2out_0 enable_0/and_2/a_n26_14# vdd enable_0/and_2/w_26_9# CMOSP w=7 l=4
+  ad=184 pd=80 as=0 ps=0
M1031 vdd a2 enable_0/and_2/a_n26_14# enable_0/and_2/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1032 a2out_0 enable_0/and_2/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=309 pd=102 as=0 ps=0
M1033 enable_0/and_2/a_n26_14# enable_0/en vdd enable_0/and_2/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1034 enable_0/and_2/a_n26_n23# enable_0/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1035 enable_0/and_2/a_n26_14# a2 enable_0/and_2/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1036 a3out_0 enable_0/and_3/a_n26_14# vdd enable_0/and_3/w_26_9# CMOSP w=7 l=4
+  ad=184 pd=80 as=0 ps=0
M1037 vdd a3 enable_0/and_3/a_n26_14# enable_0/and_3/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1038 a3out_0 enable_0/and_3/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=309 pd=102 as=0 ps=0
M1039 enable_0/and_3/a_n26_14# enable_0/en vdd enable_0/and_3/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1040 enable_0/and_3/a_n26_n23# enable_0/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1041 enable_0/and_3/a_n26_14# a3 enable_0/and_3/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1042 b0out_0 enable_0/and_4/a_n26_14# vdd enable_0/and_4/w_26_9# CMOSP w=7 l=4
+  ad=184 pd=80 as=0 ps=0
M1043 vdd b0 enable_0/and_4/a_n26_14# enable_0/and_4/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1044 b0out_0 enable_0/and_4/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=309 pd=102 as=0 ps=0
M1045 enable_0/and_4/a_n26_14# enable_0/en vdd enable_0/and_4/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1046 enable_0/and_4/a_n26_n23# enable_0/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1047 enable_0/and_4/a_n26_14# b0 enable_0/and_4/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1048 b1out_1 enable_1/and_5/a_n26_14# vdd enable_1/and_5/w_26_9# CMOSP w=7 l=4
+  ad=184 pd=80 as=0 ps=0
M1049 vdd b1 enable_1/and_5/a_n26_14# enable_1/and_5/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1050 b1out_1 enable_1/and_5/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=309 pd=102 as=0 ps=0
M1051 enable_1/and_5/a_n26_14# enable_1/en vdd enable_1/and_5/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1052 enable_1/and_5/a_n26_n23# enable_1/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1053 enable_1/and_5/a_n26_14# b1 enable_1/and_5/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1054 b3out_1 enable_1/and_7/a_n26_14# vdd enable_1/and_7/w_26_9# CMOSP w=7 l=4
+  ad=184 pd=80 as=0 ps=0
M1055 vdd b3 enable_1/and_7/a_n26_14# enable_1/and_7/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1056 b3out_1 enable_1/and_7/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=309 pd=102 as=0 ps=0
M1057 enable_1/and_7/a_n26_14# enable_1/en vdd enable_1/and_7/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1058 enable_1/and_7/a_n26_n23# enable_1/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1059 enable_1/and_7/a_n26_14# b3 enable_1/and_7/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1060 b2out_1 enable_1/and_6/a_n26_14# vdd enable_1/and_6/w_26_9# CMOSP w=7 l=4
+  ad=184 pd=80 as=0 ps=0
M1061 vdd b2 enable_1/and_6/a_n26_14# enable_1/and_6/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1062 b2out_1 enable_1/and_6/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=309 pd=102 as=0 ps=0
M1063 enable_1/and_6/a_n26_14# enable_1/en vdd enable_1/and_6/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1064 enable_1/and_6/a_n26_n23# enable_1/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1065 enable_1/and_6/a_n26_14# b2 enable_1/and_6/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1066 a0_out1 enable_1/and_0/a_n26_14# vdd enable_1/and_0/w_26_9# CMOSP w=7 l=4
+  ad=184 pd=80 as=0 ps=0
M1067 vdd a0 enable_1/and_0/a_n26_14# enable_1/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1068 a0_out1 enable_1/and_0/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=309 pd=102 as=0 ps=0
M1069 enable_1/and_0/a_n26_14# enable_1/en vdd enable_1/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1070 enable_1/and_0/a_n26_n23# enable_1/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1071 enable_1/and_0/a_n26_14# a0 enable_1/and_0/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1072 a1out_1 enable_1/and_1/a_n26_14# vdd enable_1/and_1/w_26_9# CMOSP w=7 l=4
+  ad=184 pd=80 as=0 ps=0
M1073 vdd a1 enable_1/and_1/a_n26_14# enable_1/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1074 a1out_1 enable_1/and_1/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=309 pd=102 as=0 ps=0
M1075 enable_1/and_1/a_n26_14# enable_1/en vdd enable_1/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1076 enable_1/and_1/a_n26_n23# enable_1/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1077 enable_1/and_1/a_n26_14# a1 enable_1/and_1/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1078 a2out_1 enable_1/and_2/a_n26_14# vdd enable_1/and_2/w_26_9# CMOSP w=7 l=4
+  ad=184 pd=80 as=0 ps=0
M1079 vdd a2 enable_1/and_2/a_n26_14# enable_1/and_2/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1080 a2out_1 enable_1/and_2/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=309 pd=102 as=0 ps=0
M1081 enable_1/and_2/a_n26_14# enable_1/en vdd enable_1/and_2/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1082 enable_1/and_2/a_n26_n23# enable_1/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1083 enable_1/and_2/a_n26_14# a2 enable_1/and_2/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1084 a3out_1 enable_1/and_3/a_n26_14# vdd enable_1/and_3/w_26_9# CMOSP w=7 l=4
+  ad=184 pd=80 as=0 ps=0
M1085 vdd a3 enable_1/and_3/a_n26_14# enable_1/and_3/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1086 a3out_1 enable_1/and_3/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=309 pd=102 as=0 ps=0
M1087 enable_1/and_3/a_n26_14# enable_1/en vdd enable_1/and_3/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1088 enable_1/and_3/a_n26_n23# enable_1/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1089 enable_1/and_3/a_n26_14# a3 enable_1/and_3/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1090 b0out_1 enable_1/and_4/a_n26_14# vdd enable_1/and_4/w_26_9# CMOSP w=7 l=4
+  ad=184 pd=80 as=0 ps=0
M1091 vdd b0 enable_1/and_4/a_n26_14# enable_1/and_4/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1092 b0out_1 enable_1/and_4/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=309 pd=102 as=0 ps=0
M1093 enable_1/and_4/a_n26_14# enable_1/en vdd enable_1/and_4/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1094 enable_1/and_4/a_n26_n23# enable_1/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1095 enable_1/and_4/a_n26_14# b0 enable_1/and_4/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1096 b1out_2 enable_2/and_5/a_n26_14# vdd enable_2/and_5/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1097 vdd b1 enable_2/and_5/a_n26_14# enable_2/and_5/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1098 b1out_2 enable_2/and_5/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1099 enable_2/and_5/a_n26_14# enable_2/en vdd enable_2/and_5/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1100 enable_2/and_5/a_n26_n23# enable_2/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1101 enable_2/and_5/a_n26_14# b1 enable_2/and_5/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1102 b3out_2 enable_2/and_7/a_n26_14# vdd enable_2/and_7/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1103 vdd b3 enable_2/and_7/a_n26_14# enable_2/and_7/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1104 b3out_2 enable_2/and_7/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1105 enable_2/and_7/a_n26_14# enable_2/en vdd enable_2/and_7/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1106 enable_2/and_7/a_n26_n23# enable_2/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1107 enable_2/and_7/a_n26_14# b3 enable_2/and_7/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1108 b2out_2 enable_2/and_6/a_n26_14# vdd enable_2/and_6/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1109 vdd b2 enable_2/and_6/a_n26_14# enable_2/and_6/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1110 b2out_2 enable_2/and_6/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1111 enable_2/and_6/a_n26_14# enable_2/en vdd enable_2/and_6/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1112 enable_2/and_6/a_n26_n23# enable_2/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1113 enable_2/and_6/a_n26_14# b2 enable_2/and_6/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1114 a0out_2 enable_2/and_0/a_n26_14# vdd enable_2/and_0/w_26_9# CMOSP w=7 l=4
+  ad=184 pd=80 as=0 ps=0
M1115 vdd a0 enable_2/and_0/a_n26_14# enable_2/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1116 a0out_2 enable_2/and_0/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=309 pd=102 as=0 ps=0
M1117 enable_2/and_0/a_n26_14# enable_2/en vdd enable_2/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1118 enable_2/and_0/a_n26_n23# enable_2/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1119 enable_2/and_0/a_n26_14# a0 enable_2/and_0/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1120 a1out_2 enable_2/and_1/a_n26_14# vdd enable_2/and_1/w_26_9# CMOSP w=7 l=4
+  ad=184 pd=80 as=0 ps=0
M1121 vdd a1 enable_2/and_1/a_n26_14# enable_2/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1122 a1out_2 enable_2/and_1/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=309 pd=102 as=0 ps=0
M1123 enable_2/and_1/a_n26_14# enable_2/en vdd enable_2/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1124 enable_2/and_1/a_n26_n23# enable_2/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1125 enable_2/and_1/a_n26_14# a1 enable_2/and_1/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1126 a2out_2 enable_2/and_2/a_n26_14# vdd enable_2/and_2/w_26_9# CMOSP w=7 l=4
+  ad=184 pd=80 as=0 ps=0
M1127 vdd a2 enable_2/and_2/a_n26_14# enable_2/and_2/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1128 a2out_2 enable_2/and_2/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=309 pd=102 as=0 ps=0
M1129 enable_2/and_2/a_n26_14# enable_2/en vdd enable_2/and_2/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1130 enable_2/and_2/a_n26_n23# enable_2/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1131 enable_2/and_2/a_n26_14# a2 enable_2/and_2/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1132 a3out_2 enable_2/and_3/a_n26_14# vdd enable_2/and_3/w_26_9# CMOSP w=7 l=4
+  ad=184 pd=80 as=0 ps=0
M1133 vdd a3 enable_2/and_3/a_n26_14# enable_2/and_3/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1134 a3out_2 enable_2/and_3/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=309 pd=102 as=0 ps=0
M1135 enable_2/and_3/a_n26_14# enable_2/en vdd enable_2/and_3/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1136 enable_2/and_3/a_n26_n23# enable_2/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1137 enable_2/and_3/a_n26_14# a3 enable_2/and_3/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1138 boout_2 enable_2/and_4/a_n26_14# vdd enable_2/and_4/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1139 vdd b0 enable_2/and_4/a_n26_14# enable_2/and_4/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1140 boout_2 enable_2/and_4/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1141 enable_2/and_4/a_n26_14# enable_2/en vdd enable_2/and_4/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1142 enable_2/and_4/a_n26_n23# enable_2/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1143 enable_2/and_4/a_n26_14# b0 enable_2/and_4/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1144 b1out_3 enable_3/and_5/a_n26_14# vdd enable_3/and_5/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1145 vdd b1 enable_3/and_5/a_n26_14# enable_3/and_5/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1146 b1out_3 enable_3/and_5/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1147 enable_3/and_5/a_n26_14# enable_3/en vdd enable_3/and_5/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1148 enable_3/and_5/a_n26_n23# enable_3/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1149 enable_3/and_5/a_n26_14# b1 enable_3/and_5/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1150 b3out_3 enable_3/and_7/a_n26_14# vdd enable_3/and_7/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1151 vdd b3 enable_3/and_7/a_n26_14# enable_3/and_7/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1152 b3out_3 enable_3/and_7/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1153 enable_3/and_7/a_n26_14# enable_3/en vdd enable_3/and_7/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1154 enable_3/and_7/a_n26_n23# enable_3/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1155 enable_3/and_7/a_n26_14# b3 enable_3/and_7/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1156 b2out_3 enable_3/and_6/a_n26_14# vdd enable_3/and_6/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1157 vdd b2 enable_3/and_6/a_n26_14# enable_3/and_6/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1158 b2out_3 enable_3/and_6/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1159 enable_3/and_6/a_n26_14# enable_3/en vdd enable_3/and_6/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1160 enable_3/and_6/a_n26_n23# enable_3/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1161 enable_3/and_6/a_n26_14# b2 enable_3/and_6/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1162 a0out_3 enable_3/and_0/a_n26_14# vdd enable_3/and_0/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1163 vdd a0 enable_3/and_0/a_n26_14# enable_3/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1164 a0out_3 enable_3/and_0/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1165 enable_3/and_0/a_n26_14# enable_3/en vdd enable_3/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1166 enable_3/and_0/a_n26_n23# enable_3/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1167 enable_3/and_0/a_n26_14# a0 enable_3/and_0/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1168 a1out_3 enable_3/and_1/a_n26_14# vdd enable_3/and_1/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1169 vdd a1 enable_3/and_1/a_n26_14# enable_3/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1170 a1out_3 enable_3/and_1/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1171 enable_3/and_1/a_n26_14# enable_3/en vdd enable_3/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1172 enable_3/and_1/a_n26_n23# enable_3/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1173 enable_3/and_1/a_n26_14# a1 enable_3/and_1/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1174 a2out_3 enable_3/and_2/a_n26_14# vdd enable_3/and_2/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1175 vdd a2 enable_3/and_2/a_n26_14# enable_3/and_2/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1176 a2out_3 enable_3/and_2/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1177 enable_3/and_2/a_n26_14# enable_3/en vdd enable_3/and_2/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1178 enable_3/and_2/a_n26_n23# enable_3/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1179 enable_3/and_2/a_n26_14# a2 enable_3/and_2/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1180 a3out_3 enable_3/and_3/a_n26_14# vdd enable_3/and_3/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1181 vdd a3 enable_3/and_3/a_n26_14# enable_3/and_3/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1182 a3out_3 enable_3/and_3/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1183 enable_3/and_3/a_n26_14# enable_3/en vdd enable_3/and_3/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1184 enable_3/and_3/a_n26_n23# enable_3/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1185 enable_3/and_3/a_n26_14# a3 enable_3/and_3/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1186 b0out_3 enable_3/and_4/a_n26_14# vdd enable_3/and_4/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1187 vdd b0 enable_3/and_4/a_n26_14# enable_3/and_4/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1188 b0out_3 enable_3/and_4/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1189 enable_3/and_4/a_n26_14# enable_3/en vdd enable_3/and_4/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1190 enable_3/and_4/a_n26_n23# enable_3/en gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1191 enable_3/and_4/a_n26_14# b0 enable_3/and_4/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1192 out0 AND_Block_0/and_0/a_n26_14# vdd AND_Block_0/and_0/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1193 vdd b0out_3 AND_Block_0/and_0/a_n26_14# AND_Block_0/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1194 out0 AND_Block_0/and_0/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1195 AND_Block_0/and_0/a_n26_14# a0out_3 vdd AND_Block_0/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1196 AND_Block_0/and_0/a_n26_n23# a0out_3 gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1197 AND_Block_0/and_0/a_n26_14# b0out_3 AND_Block_0/and_0/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1198 out1 AND_Block_0/and_1/a_n26_14# vdd AND_Block_0/and_1/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1199 vdd b1out_3 AND_Block_0/and_1/a_n26_14# AND_Block_0/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1200 out1 AND_Block_0/and_1/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1201 AND_Block_0/and_1/a_n26_14# a1out_3 vdd AND_Block_0/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1202 AND_Block_0/and_1/a_n26_n23# a1out_3 gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1203 AND_Block_0/and_1/a_n26_14# b1out_3 AND_Block_0/and_1/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1204 out2 AND_Block_0/and_2/a_n26_14# vdd AND_Block_0/and_2/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1205 vdd b2out_3 AND_Block_0/and_2/a_n26_14# AND_Block_0/and_2/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1206 out2 AND_Block_0/and_2/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1207 AND_Block_0/and_2/a_n26_14# a2out_3 vdd AND_Block_0/and_2/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1208 AND_Block_0/and_2/a_n26_n23# a2out_3 gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1209 AND_Block_0/and_2/a_n26_14# b2out_3 AND_Block_0/and_2/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1210 out3 AND_Block_0/and_3/a_n26_14# vdd AND_Block_0/and_3/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1211 vdd b3out_3 AND_Block_0/and_3/a_n26_14# AND_Block_0/and_3/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1212 out3 AND_Block_0/and_3/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1213 AND_Block_0/and_3/a_n26_14# a3out_3 vdd AND_Block_0/and_3/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1214 AND_Block_0/and_3/a_n26_n23# a3out_3 gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1215 AND_Block_0/and_3/a_n26_14# b3out_3 AND_Block_0/and_3/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1216 4bitadder_0/fulladder_0/or_0/a_n15_32# 4bitadder_0/fulladder_0/or_0/a gnd Gnd CMOSN w=16 l=5
+  ad=304 pd=70 as=0 ps=0
M1217 4bitadder_0/c1 4bitadder_0/fulladder_0/or_0/a_n15_32# vdd 4bitadder_0/fulladder_0/or_0/w_58_101# CMOSP w=16 l=6
+  ad=288 pd=68 as=0 ps=0
M1218 gnd 4bitadder_0/fulladder_0/or_0/b 4bitadder_0/fulladder_0/or_0/a_n15_32# Gnd CMOSN w=16 l=5
+  ad=0 pd=0 as=0 ps=0
M1219 4bitadder_0/fulladder_0/or_0/a_n15_32# 4bitadder_0/fulladder_0/or_0/b 4bitadder_0/fulladder_0/or_0/a_n15_107# 4bitadder_0/fulladder_0/or_0/w_n48_101# CMOSP w=16 l=5
+  ad=448 pd=88 as=304 ps=70
M1220 4bitadder_0/c1 4bitadder_0/fulladder_0/or_0/a_n15_32# gnd Gnd CMOSN w=16 l=6
+  ad=320 pd=72 as=0 ps=0
M1221 4bitadder_0/fulladder_0/or_0/a_n15_107# 4bitadder_0/fulladder_0/or_0/a vdd 4bitadder_0/fulladder_0/or_0/w_n48_101# CMOSP w=16 l=5
+  ad=0 pd=0 as=0 ps=0
M1222 4bitadder_0/fulladder_0/or_0/a 4bitadder_0/fulladder_0/and_0/a_n26_14# vdd 4bitadder_0/fulladder_0/and_0/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1223 vdd s0 4bitadder_0/fulladder_0/and_0/a_n26_14# 4bitadder_0/fulladder_0/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1224 4bitadder_0/fulladder_0/or_0/a 4bitadder_0/fulladder_0/and_0/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1225 4bitadder_0/fulladder_0/and_0/a_n26_14# 4bitadder_0/fulladder_0/axorb vdd 4bitadder_0/fulladder_0/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1226 4bitadder_0/fulladder_0/and_0/a_n26_n23# 4bitadder_0/fulladder_0/axorb gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1227 4bitadder_0/fulladder_0/and_0/a_n26_14# s0 4bitadder_0/fulladder_0/and_0/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1228 4bitadder_0/fulladder_0/axorb 4bitadder_0/b0xorM 4bitadder_0/fulladder_0/XOR_0/abar Gnd CMOSN w=11 l=6
+  ad=495 pd=156 as=407 ps=118
M1229 4bitadder_0/fulladder_0/XOR_0/bbar 4bitadder_0/b0xorM gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1230 4bitadder_0/fulladder_0/axorb 4bitadder_0/fulladder_0/XOR_0/bbar 4bitadder_0/fulladder_0/XOR_0/abar 4bitadder_0/fulladder_0/XOR_0/w_62_n20# CMOSP w=12 l=6
+  ad=252 pd=110 as=218 ps=84
M1231 vdd 4bitadder_0/b0xorM 4bitadder_0/fulladder_0/XOR_0/bbar 4bitadder_0/fulladder_0/XOR_0/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1232 4bitadder_0/fulladder_0/axorb 4bitadder_0/b0xorM a0out_0 4bitadder_0/fulladder_0/XOR_0/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1233 4bitadder_0/fulladder_0/XOR_0/abar a0out_0 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1234 vdd a0out_0 4bitadder_0/fulladder_0/XOR_0/abar 4bitadder_0/fulladder_0/XOR_0/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1235 4bitadder_0/fulladder_0/axorb 4bitadder_0/fulladder_0/XOR_0/bbar a0out_0 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1236 4bitadder_0/fulladder_0/or_0/b 4bitadder_0/fulladder_0/and_1/a_n26_14# vdd 4bitadder_0/fulladder_0/and_1/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1237 vdd a0out_0 4bitadder_0/fulladder_0/and_1/a_n26_14# 4bitadder_0/fulladder_0/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1238 4bitadder_0/fulladder_0/or_0/b 4bitadder_0/fulladder_0/and_1/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1239 4bitadder_0/fulladder_0/and_1/a_n26_14# 4bitadder_0/b0xorM vdd 4bitadder_0/fulladder_0/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1240 4bitadder_0/fulladder_0/and_1/a_n26_n23# 4bitadder_0/b0xorM gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1241 4bitadder_0/fulladder_0/and_1/a_n26_14# a0out_0 4bitadder_0/fulladder_0/and_1/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1242 s0_add s0 4bitadder_0/fulladder_0/XOR_1/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1243 4bitadder_0/fulladder_0/XOR_1/bbar s0 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1244 s0_add 4bitadder_0/fulladder_0/XOR_1/bbar 4bitadder_0/fulladder_0/XOR_1/abar 4bitadder_0/fulladder_0/XOR_1/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1245 vdd s0 4bitadder_0/fulladder_0/XOR_1/bbar 4bitadder_0/fulladder_0/XOR_1/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1246 s0_add s0 4bitadder_0/fulladder_0/axorb 4bitadder_0/fulladder_0/XOR_1/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1247 4bitadder_0/fulladder_0/XOR_1/abar 4bitadder_0/fulladder_0/axorb gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1248 vdd 4bitadder_0/fulladder_0/axorb 4bitadder_0/fulladder_0/XOR_1/abar 4bitadder_0/fulladder_0/XOR_1/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1249 s0_add 4bitadder_0/fulladder_0/XOR_1/bbar 4bitadder_0/fulladder_0/axorb Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1250 4bitadder_0/fulladder_1/or_0/a_n15_32# 4bitadder_0/fulladder_1/or_0/a gnd Gnd CMOSN w=16 l=5
+  ad=304 pd=70 as=0 ps=0
M1251 4bitadder_0/c2 4bitadder_0/fulladder_1/or_0/a_n15_32# vdd 4bitadder_0/fulladder_1/or_0/w_58_101# CMOSP w=16 l=6
+  ad=288 pd=68 as=0 ps=0
M1252 gnd 4bitadder_0/fulladder_1/or_0/b 4bitadder_0/fulladder_1/or_0/a_n15_32# Gnd CMOSN w=16 l=5
+  ad=0 pd=0 as=0 ps=0
M1253 4bitadder_0/fulladder_1/or_0/a_n15_32# 4bitadder_0/fulladder_1/or_0/b 4bitadder_0/fulladder_1/or_0/a_n15_107# 4bitadder_0/fulladder_1/or_0/w_n48_101# CMOSP w=16 l=5
+  ad=448 pd=88 as=304 ps=70
M1254 4bitadder_0/c2 4bitadder_0/fulladder_1/or_0/a_n15_32# gnd Gnd CMOSN w=16 l=6
+  ad=320 pd=72 as=0 ps=0
M1255 4bitadder_0/fulladder_1/or_0/a_n15_107# 4bitadder_0/fulladder_1/or_0/a vdd 4bitadder_0/fulladder_1/or_0/w_n48_101# CMOSP w=16 l=5
+  ad=0 pd=0 as=0 ps=0
M1256 4bitadder_0/fulladder_1/or_0/a 4bitadder_0/fulladder_1/and_0/a_n26_14# vdd 4bitadder_0/fulladder_1/and_0/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1257 vdd 4bitadder_0/c1 4bitadder_0/fulladder_1/and_0/a_n26_14# 4bitadder_0/fulladder_1/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1258 4bitadder_0/fulladder_1/or_0/a 4bitadder_0/fulladder_1/and_0/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1259 4bitadder_0/fulladder_1/and_0/a_n26_14# 4bitadder_0/fulladder_1/axorb vdd 4bitadder_0/fulladder_1/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1260 4bitadder_0/fulladder_1/and_0/a_n26_n23# 4bitadder_0/fulladder_1/axorb gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1261 4bitadder_0/fulladder_1/and_0/a_n26_14# 4bitadder_0/c1 4bitadder_0/fulladder_1/and_0/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1262 4bitadder_0/fulladder_1/axorb 4bitadder_0/XOR_1/out 4bitadder_0/fulladder_1/XOR_0/abar Gnd CMOSN w=11 l=6
+  ad=495 pd=156 as=407 ps=118
M1263 4bitadder_0/fulladder_1/XOR_0/bbar 4bitadder_0/XOR_1/out gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1264 4bitadder_0/fulladder_1/axorb 4bitadder_0/fulladder_1/XOR_0/bbar 4bitadder_0/fulladder_1/XOR_0/abar 4bitadder_0/fulladder_1/XOR_0/w_62_n20# CMOSP w=12 l=6
+  ad=252 pd=110 as=218 ps=84
M1265 vdd 4bitadder_0/XOR_1/out 4bitadder_0/fulladder_1/XOR_0/bbar 4bitadder_0/fulladder_1/XOR_0/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1266 4bitadder_0/fulladder_1/axorb 4bitadder_0/XOR_1/out a1out_0 4bitadder_0/fulladder_1/XOR_0/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1267 4bitadder_0/fulladder_1/XOR_0/abar a1out_0 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1268 vdd a1out_0 4bitadder_0/fulladder_1/XOR_0/abar 4bitadder_0/fulladder_1/XOR_0/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1269 4bitadder_0/fulladder_1/axorb 4bitadder_0/fulladder_1/XOR_0/bbar a1out_0 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1270 4bitadder_0/fulladder_1/or_0/b 4bitadder_0/fulladder_1/and_1/a_n26_14# vdd 4bitadder_0/fulladder_1/and_1/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1271 vdd a1out_0 4bitadder_0/fulladder_1/and_1/a_n26_14# 4bitadder_0/fulladder_1/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1272 4bitadder_0/fulladder_1/or_0/b 4bitadder_0/fulladder_1/and_1/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1273 4bitadder_0/fulladder_1/and_1/a_n26_14# 4bitadder_0/XOR_1/out vdd 4bitadder_0/fulladder_1/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1274 4bitadder_0/fulladder_1/and_1/a_n26_n23# 4bitadder_0/XOR_1/out gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1275 4bitadder_0/fulladder_1/and_1/a_n26_14# a1out_0 4bitadder_0/fulladder_1/and_1/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1276 s1_add 4bitadder_0/c1 4bitadder_0/fulladder_1/XOR_1/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1277 4bitadder_0/fulladder_1/XOR_1/bbar 4bitadder_0/c1 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1278 s1_add 4bitadder_0/fulladder_1/XOR_1/bbar 4bitadder_0/fulladder_1/XOR_1/abar 4bitadder_0/fulladder_1/XOR_1/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1279 vdd 4bitadder_0/c1 4bitadder_0/fulladder_1/XOR_1/bbar 4bitadder_0/fulladder_1/XOR_1/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1280 s1_add 4bitadder_0/c1 4bitadder_0/fulladder_1/axorb 4bitadder_0/fulladder_1/XOR_1/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1281 4bitadder_0/fulladder_1/XOR_1/abar 4bitadder_0/fulladder_1/axorb gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1282 vdd 4bitadder_0/fulladder_1/axorb 4bitadder_0/fulladder_1/XOR_1/abar 4bitadder_0/fulladder_1/XOR_1/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1283 s1_add 4bitadder_0/fulladder_1/XOR_1/bbar 4bitadder_0/fulladder_1/axorb Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1284 4bitadder_0/fulladder_2/or_0/a_n15_32# 4bitadder_0/fulladder_2/or_0/a gnd Gnd CMOSN w=16 l=5
+  ad=304 pd=70 as=0 ps=0
M1285 4bitadder_0/c3 4bitadder_0/fulladder_2/or_0/a_n15_32# vdd 4bitadder_0/fulladder_2/or_0/w_58_101# CMOSP w=16 l=6
+  ad=288 pd=68 as=0 ps=0
M1286 gnd 4bitadder_0/fulladder_2/or_0/b 4bitadder_0/fulladder_2/or_0/a_n15_32# Gnd CMOSN w=16 l=5
+  ad=0 pd=0 as=0 ps=0
M1287 4bitadder_0/fulladder_2/or_0/a_n15_32# 4bitadder_0/fulladder_2/or_0/b 4bitadder_0/fulladder_2/or_0/a_n15_107# 4bitadder_0/fulladder_2/or_0/w_n48_101# CMOSP w=16 l=5
+  ad=448 pd=88 as=304 ps=70
M1288 4bitadder_0/c3 4bitadder_0/fulladder_2/or_0/a_n15_32# gnd Gnd CMOSN w=16 l=6
+  ad=320 pd=72 as=0 ps=0
M1289 4bitadder_0/fulladder_2/or_0/a_n15_107# 4bitadder_0/fulladder_2/or_0/a vdd 4bitadder_0/fulladder_2/or_0/w_n48_101# CMOSP w=16 l=5
+  ad=0 pd=0 as=0 ps=0
M1290 4bitadder_0/fulladder_2/or_0/a 4bitadder_0/fulladder_2/and_0/a_n26_14# vdd 4bitadder_0/fulladder_2/and_0/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1291 vdd 4bitadder_0/c2 4bitadder_0/fulladder_2/and_0/a_n26_14# 4bitadder_0/fulladder_2/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1292 4bitadder_0/fulladder_2/or_0/a 4bitadder_0/fulladder_2/and_0/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1293 4bitadder_0/fulladder_2/and_0/a_n26_14# 4bitadder_0/fulladder_2/axorb vdd 4bitadder_0/fulladder_2/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1294 4bitadder_0/fulladder_2/and_0/a_n26_n23# 4bitadder_0/fulladder_2/axorb gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1295 4bitadder_0/fulladder_2/and_0/a_n26_14# 4bitadder_0/c2 4bitadder_0/fulladder_2/and_0/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1296 4bitadder_0/fulladder_2/axorb 4bitadder_0/XOR_2/out 4bitadder_0/fulladder_2/XOR_0/abar Gnd CMOSN w=11 l=6
+  ad=495 pd=156 as=407 ps=118
M1297 4bitadder_0/fulladder_2/XOR_0/bbar 4bitadder_0/XOR_2/out gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1298 4bitadder_0/fulladder_2/axorb 4bitadder_0/fulladder_2/XOR_0/bbar 4bitadder_0/fulladder_2/XOR_0/abar 4bitadder_0/fulladder_2/XOR_0/w_62_n20# CMOSP w=12 l=6
+  ad=252 pd=110 as=218 ps=84
M1299 vdd 4bitadder_0/XOR_2/out 4bitadder_0/fulladder_2/XOR_0/bbar 4bitadder_0/fulladder_2/XOR_0/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1300 4bitadder_0/fulladder_2/axorb 4bitadder_0/XOR_2/out a2out_0 4bitadder_0/fulladder_2/XOR_0/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1301 4bitadder_0/fulladder_2/XOR_0/abar a2out_0 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1302 vdd a2out_0 4bitadder_0/fulladder_2/XOR_0/abar 4bitadder_0/fulladder_2/XOR_0/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1303 4bitadder_0/fulladder_2/axorb 4bitadder_0/fulladder_2/XOR_0/bbar a2out_0 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1304 4bitadder_0/fulladder_2/or_0/b 4bitadder_0/fulladder_2/and_1/a_n26_14# vdd 4bitadder_0/fulladder_2/and_1/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1305 vdd a2out_0 4bitadder_0/fulladder_2/and_1/a_n26_14# 4bitadder_0/fulladder_2/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1306 4bitadder_0/fulladder_2/or_0/b 4bitadder_0/fulladder_2/and_1/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1307 4bitadder_0/fulladder_2/and_1/a_n26_14# 4bitadder_0/XOR_2/out vdd 4bitadder_0/fulladder_2/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1308 4bitadder_0/fulladder_2/and_1/a_n26_n23# 4bitadder_0/XOR_2/out gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1309 4bitadder_0/fulladder_2/and_1/a_n26_14# a2out_0 4bitadder_0/fulladder_2/and_1/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1310 s2_add 4bitadder_0/c2 4bitadder_0/fulladder_2/XOR_1/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1311 4bitadder_0/fulladder_2/XOR_1/bbar 4bitadder_0/c2 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1312 s2_add 4bitadder_0/fulladder_2/XOR_1/bbar 4bitadder_0/fulladder_2/XOR_1/abar 4bitadder_0/fulladder_2/XOR_1/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1313 vdd 4bitadder_0/c2 4bitadder_0/fulladder_2/XOR_1/bbar 4bitadder_0/fulladder_2/XOR_1/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1314 s2_add 4bitadder_0/c2 4bitadder_0/fulladder_2/axorb 4bitadder_0/fulladder_2/XOR_1/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1315 4bitadder_0/fulladder_2/XOR_1/abar 4bitadder_0/fulladder_2/axorb gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1316 vdd 4bitadder_0/fulladder_2/axorb 4bitadder_0/fulladder_2/XOR_1/abar 4bitadder_0/fulladder_2/XOR_1/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1317 s2_add 4bitadder_0/fulladder_2/XOR_1/bbar 4bitadder_0/fulladder_2/axorb Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1318 4bitadder_0/fulladder_3/or_0/a_n15_32# 4bitadder_0/fulladder_3/or_0/a gnd Gnd CMOSN w=16 l=5
+  ad=304 pd=70 as=0 ps=0
M1319 fc_add 4bitadder_0/fulladder_3/or_0/a_n15_32# vdd 4bitadder_0/fulladder_3/or_0/w_58_101# CMOSP w=16 l=6
+  ad=288 pd=68 as=0 ps=0
M1320 gnd 4bitadder_0/fulladder_3/or_0/b 4bitadder_0/fulladder_3/or_0/a_n15_32# Gnd CMOSN w=16 l=5
+  ad=0 pd=0 as=0 ps=0
M1321 4bitadder_0/fulladder_3/or_0/a_n15_32# 4bitadder_0/fulladder_3/or_0/b 4bitadder_0/fulladder_3/or_0/a_n15_107# 4bitadder_0/fulladder_3/or_0/w_n48_101# CMOSP w=16 l=5
+  ad=448 pd=88 as=304 ps=70
M1322 fc_add 4bitadder_0/fulladder_3/or_0/a_n15_32# gnd Gnd CMOSN w=16 l=6
+  ad=320 pd=72 as=0 ps=0
M1323 4bitadder_0/fulladder_3/or_0/a_n15_107# 4bitadder_0/fulladder_3/or_0/a vdd 4bitadder_0/fulladder_3/or_0/w_n48_101# CMOSP w=16 l=5
+  ad=0 pd=0 as=0 ps=0
M1324 4bitadder_0/fulladder_3/or_0/a 4bitadder_0/fulladder_3/and_0/a_n26_14# vdd 4bitadder_0/fulladder_3/and_0/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1325 vdd 4bitadder_0/c3 4bitadder_0/fulladder_3/and_0/a_n26_14# 4bitadder_0/fulladder_3/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1326 4bitadder_0/fulladder_3/or_0/a 4bitadder_0/fulladder_3/and_0/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1327 4bitadder_0/fulladder_3/and_0/a_n26_14# 4bitadder_0/fulladder_3/axorb vdd 4bitadder_0/fulladder_3/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1328 4bitadder_0/fulladder_3/and_0/a_n26_n23# 4bitadder_0/fulladder_3/axorb gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1329 4bitadder_0/fulladder_3/and_0/a_n26_14# 4bitadder_0/c3 4bitadder_0/fulladder_3/and_0/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1330 4bitadder_0/fulladder_3/axorb 4bitadder_0/XOR_3/out 4bitadder_0/fulladder_3/XOR_0/abar Gnd CMOSN w=11 l=6
+  ad=495 pd=156 as=407 ps=118
M1331 4bitadder_0/fulladder_3/XOR_0/bbar 4bitadder_0/XOR_3/out gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1332 4bitadder_0/fulladder_3/axorb 4bitadder_0/fulladder_3/XOR_0/bbar 4bitadder_0/fulladder_3/XOR_0/abar 4bitadder_0/fulladder_3/XOR_0/w_62_n20# CMOSP w=12 l=6
+  ad=252 pd=110 as=218 ps=84
M1333 vdd 4bitadder_0/XOR_3/out 4bitadder_0/fulladder_3/XOR_0/bbar 4bitadder_0/fulladder_3/XOR_0/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1334 4bitadder_0/fulladder_3/axorb 4bitadder_0/XOR_3/out a3out_0 4bitadder_0/fulladder_3/XOR_0/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1335 4bitadder_0/fulladder_3/XOR_0/abar a3out_0 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1336 vdd a3out_0 4bitadder_0/fulladder_3/XOR_0/abar 4bitadder_0/fulladder_3/XOR_0/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1337 4bitadder_0/fulladder_3/axorb 4bitadder_0/fulladder_3/XOR_0/bbar a3out_0 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1338 4bitadder_0/fulladder_3/or_0/b 4bitadder_0/fulladder_3/and_1/a_n26_14# vdd 4bitadder_0/fulladder_3/and_1/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1339 vdd a3out_0 4bitadder_0/fulladder_3/and_1/a_n26_14# 4bitadder_0/fulladder_3/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1340 4bitadder_0/fulladder_3/or_0/b 4bitadder_0/fulladder_3/and_1/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1341 4bitadder_0/fulladder_3/and_1/a_n26_14# 4bitadder_0/XOR_3/out vdd 4bitadder_0/fulladder_3/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1342 4bitadder_0/fulladder_3/and_1/a_n26_n23# 4bitadder_0/XOR_3/out gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1343 4bitadder_0/fulladder_3/and_1/a_n26_14# a3out_0 4bitadder_0/fulladder_3/and_1/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1344 s3_add 4bitadder_0/c3 4bitadder_0/fulladder_3/XOR_1/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1345 4bitadder_0/fulladder_3/XOR_1/bbar 4bitadder_0/c3 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1346 s3_add 4bitadder_0/fulladder_3/XOR_1/bbar 4bitadder_0/fulladder_3/XOR_1/abar 4bitadder_0/fulladder_3/XOR_1/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1347 vdd 4bitadder_0/c3 4bitadder_0/fulladder_3/XOR_1/bbar 4bitadder_0/fulladder_3/XOR_1/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1348 s3_add 4bitadder_0/c3 4bitadder_0/fulladder_3/axorb 4bitadder_0/fulladder_3/XOR_1/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1349 4bitadder_0/fulladder_3/XOR_1/abar 4bitadder_0/fulladder_3/axorb gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1350 vdd 4bitadder_0/fulladder_3/axorb 4bitadder_0/fulladder_3/XOR_1/abar 4bitadder_0/fulladder_3/XOR_1/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1351 s3_add 4bitadder_0/fulladder_3/XOR_1/bbar 4bitadder_0/fulladder_3/axorb Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1352 4bitadder_0/b0xorM s0 4bitadder_0/XOR_0/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1353 4bitadder_0/XOR_0/bbar s0 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1354 4bitadder_0/b0xorM 4bitadder_0/XOR_0/bbar 4bitadder_0/XOR_0/abar 4bitadder_0/XOR_0/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1355 vdd s0 4bitadder_0/XOR_0/bbar 4bitadder_0/XOR_0/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1356 4bitadder_0/b0xorM s0 b0out_0 4bitadder_0/XOR_0/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1357 4bitadder_0/XOR_0/abar b0out_0 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1358 vdd b0out_0 4bitadder_0/XOR_0/abar 4bitadder_0/XOR_0/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1359 4bitadder_0/b0xorM 4bitadder_0/XOR_0/bbar b0out_0 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1360 4bitadder_0/XOR_1/out s0 4bitadder_0/XOR_1/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1361 4bitadder_0/XOR_1/bbar s0 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1362 4bitadder_0/XOR_1/out 4bitadder_0/XOR_1/bbar 4bitadder_0/XOR_1/abar 4bitadder_0/XOR_1/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1363 vdd s0 4bitadder_0/XOR_1/bbar 4bitadder_0/XOR_1/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1364 4bitadder_0/XOR_1/out s0 b1out_0 4bitadder_0/XOR_1/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1365 4bitadder_0/XOR_1/abar b1out_0 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1366 vdd b1out_0 4bitadder_0/XOR_1/abar 4bitadder_0/XOR_1/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1367 4bitadder_0/XOR_1/out 4bitadder_0/XOR_1/bbar b1out_0 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1368 4bitadder_0/XOR_2/out s0 4bitadder_0/XOR_2/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1369 4bitadder_0/XOR_2/bbar s0 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1370 4bitadder_0/XOR_2/out 4bitadder_0/XOR_2/bbar 4bitadder_0/XOR_2/abar 4bitadder_0/XOR_2/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1371 vdd s0 4bitadder_0/XOR_2/bbar 4bitadder_0/XOR_2/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1372 4bitadder_0/XOR_2/out s0 b2out_0 4bitadder_0/XOR_2/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1373 4bitadder_0/XOR_2/abar b2out_0 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1374 vdd b2out_0 4bitadder_0/XOR_2/abar 4bitadder_0/XOR_2/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1375 4bitadder_0/XOR_2/out 4bitadder_0/XOR_2/bbar b2out_0 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1376 4bitadder_0/XOR_3/out s0 4bitadder_0/XOR_3/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1377 4bitadder_0/XOR_3/bbar s0 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1378 4bitadder_0/XOR_3/out 4bitadder_0/XOR_3/bbar 4bitadder_0/XOR_3/abar 4bitadder_0/XOR_3/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1379 vdd s0 4bitadder_0/XOR_3/bbar 4bitadder_0/XOR_3/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1380 4bitadder_0/XOR_3/out s0 b3out_0 4bitadder_0/XOR_3/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1381 4bitadder_0/XOR_3/abar b3out_0 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1382 vdd b3out_0 4bitadder_0/XOR_3/abar 4bitadder_0/XOR_3/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1383 4bitadder_0/XOR_3/out 4bitadder_0/XOR_3/bbar b3out_0 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1384 comparator_0/b0bar boout_2 vdd comparator_0/not_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1385 comparator_0/b0bar boout_2 gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1386 comparator_0/b1bar b1out_2 vdd comparator_0/not_1/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1387 comparator_0/b1bar b1out_2 gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1388 agb comparator_0/4input_OR_0/y vdd comparator_0/4input_OR_0/NOT_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1389 agb comparator_0/4input_OR_0/y gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1390 vdd comparator_0/t8 comparator_0/4input_OR_0/a_n52_24# comparator_0/4input_OR_0/w_n58_n43# CMOSP w=14 l=5
+  ad=0 pd=0 as=126 ps=46
M1391 comparator_0/4input_OR_0/y comparator_0/t8 gnd Gnd CMOSN w=16 l=7
+  ad=704 pd=216 as=0 ps=0
M1392 comparator_0/4input_OR_0/a_n52_4# comparator_0/t6 comparator_0/4input_OR_0/a_n52_n15# comparator_0/4input_OR_0/w_n58_n43# CMOSP w=14 l=5
+  ad=210 pd=58 as=196 ps=56
M1393 comparator_0/4input_OR_0/y comparator_0/t5 gnd Gnd CMOSN w=16 l=7
+  ad=0 pd=0 as=0 ps=0
M1394 comparator_0/4input_OR_0/y comparator_0/t7 gnd Gnd CMOSN w=16 l=7
+  ad=0 pd=0 as=0 ps=0
M1395 comparator_0/4input_OR_0/a_n52_24# comparator_0/t7 comparator_0/4input_OR_0/a_n52_4# comparator_0/4input_OR_0/w_n58_n43# CMOSP w=14 l=5
+  ad=0 pd=0 as=0 ps=0
M1396 comparator_0/4input_OR_0/a_n52_n15# comparator_0/t5 comparator_0/4input_OR_0/y comparator_0/4input_OR_0/w_n58_n43# CMOSP w=14 l=5
+  ad=0 pd=0 as=238 ps=62
M1397 comparator_0/4input_OR_0/y comparator_0/t6 gnd Gnd CMOSN w=16 l=7
+  ad=0 pd=0 as=0 ps=0
M1398 comparator_0/b2bar b2out_2 vdd comparator_0/not_2/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1399 comparator_0/b2bar b2out_2 gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1400 comparator_0/a3xnorb3 comparator_0/xnor_0/not_0/in vdd comparator_0/xnor_0/not_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1401 comparator_0/a3xnorb3 comparator_0/xnor_0/not_0/in gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1402 comparator_0/xnor_0/not_0/in b3out_2 comparator_0/xnor_0/XOR_0/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1403 comparator_0/xnor_0/XOR_0/bbar b3out_2 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1404 comparator_0/xnor_0/not_0/in comparator_0/xnor_0/XOR_0/bbar comparator_0/xnor_0/XOR_0/abar comparator_0/xnor_0/XOR_0/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1405 vdd b3out_2 comparator_0/xnor_0/XOR_0/bbar comparator_0/xnor_0/XOR_0/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1406 comparator_0/xnor_0/not_0/in b3out_2 a3out_2 comparator_0/xnor_0/XOR_0/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1407 comparator_0/xnor_0/XOR_0/abar a3out_2 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1408 vdd a3out_2 comparator_0/xnor_0/XOR_0/abar comparator_0/xnor_0/XOR_0/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1409 comparator_0/xnor_0/not_0/in comparator_0/xnor_0/XOR_0/bbar a3out_2 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1410 comparator_0/b3bar b3out_2 vdd comparator_0/not_3/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1411 comparator_0/b3bar b3out_2 gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1412 comparator_0/a2xnorb2 comparator_0/xnor_1/not_0/in vdd comparator_0/xnor_1/not_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1413 comparator_0/a2xnorb2 comparator_0/xnor_1/not_0/in gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1414 comparator_0/xnor_1/not_0/in b2out_2 comparator_0/xnor_1/XOR_0/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1415 comparator_0/xnor_1/XOR_0/bbar b2out_2 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1416 comparator_0/xnor_1/not_0/in comparator_0/xnor_1/XOR_0/bbar comparator_0/xnor_1/XOR_0/abar comparator_0/xnor_1/XOR_0/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1417 vdd b2out_2 comparator_0/xnor_1/XOR_0/bbar comparator_0/xnor_1/XOR_0/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1418 comparator_0/xnor_1/not_0/in b2out_2 a2out_2 comparator_0/xnor_1/XOR_0/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1419 comparator_0/xnor_1/XOR_0/abar a2out_2 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1420 vdd a2out_2 comparator_0/xnor_1/XOR_0/abar comparator_0/xnor_1/XOR_0/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1421 comparator_0/xnor_1/not_0/in comparator_0/xnor_1/XOR_0/bbar a2out_2 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1422 comparator_0/a0bar a0out_2 vdd comparator_0/not_4/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1423 comparator_0/a0bar a0out_2 gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1424 bga comparator_0/4input_OR_1/y vdd comparator_0/4input_OR_1/NOT_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1425 bga comparator_0/4input_OR_1/y gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1426 vdd comparator_0/t4 comparator_0/4input_OR_1/a_n52_24# comparator_0/4input_OR_1/w_n58_n43# CMOSP w=14 l=5
+  ad=0 pd=0 as=126 ps=46
M1427 comparator_0/4input_OR_1/y comparator_0/t4 gnd Gnd CMOSN w=16 l=7
+  ad=704 pd=216 as=0 ps=0
M1428 comparator_0/4input_OR_1/a_n52_4# comparator_0/t2 comparator_0/4input_OR_1/a_n52_n15# comparator_0/4input_OR_1/w_n58_n43# CMOSP w=14 l=5
+  ad=210 pd=58 as=196 ps=56
M1429 comparator_0/4input_OR_1/y comparator_0/t1 gnd Gnd CMOSN w=16 l=7
+  ad=0 pd=0 as=0 ps=0
M1430 comparator_0/4input_OR_1/y comparator_0/t3 gnd Gnd CMOSN w=16 l=7
+  ad=0 pd=0 as=0 ps=0
M1431 comparator_0/4input_OR_1/a_n52_24# comparator_0/t3 comparator_0/4input_OR_1/a_n52_4# comparator_0/4input_OR_1/w_n58_n43# CMOSP w=14 l=5
+  ad=0 pd=0 as=0 ps=0
M1432 comparator_0/4input_OR_1/a_n52_n15# comparator_0/t1 comparator_0/4input_OR_1/y comparator_0/4input_OR_1/w_n58_n43# CMOSP w=14 l=5
+  ad=0 pd=0 as=238 ps=62
M1433 comparator_0/4input_OR_1/y comparator_0/t2 gnd Gnd CMOSN w=16 l=7
+  ad=0 pd=0 as=0 ps=0
M1434 comparator_0/a1xnorb1 comparator_0/xnor_2/not_0/in vdd comparator_0/xnor_2/not_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1435 comparator_0/a1xnorb1 comparator_0/xnor_2/not_0/in gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1436 comparator_0/xnor_2/not_0/in b1out_2 comparator_0/xnor_2/XOR_0/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1437 comparator_0/xnor_2/XOR_0/bbar b1out_2 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1438 comparator_0/xnor_2/not_0/in comparator_0/xnor_2/XOR_0/bbar comparator_0/xnor_2/XOR_0/abar comparator_0/xnor_2/XOR_0/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1439 vdd b1out_2 comparator_0/xnor_2/XOR_0/bbar comparator_0/xnor_2/XOR_0/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1440 comparator_0/xnor_2/not_0/in b1out_2 a1out_2 comparator_0/xnor_2/XOR_0/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1441 comparator_0/xnor_2/XOR_0/abar a1out_2 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1442 vdd a1out_2 comparator_0/xnor_2/XOR_0/abar comparator_0/xnor_2/XOR_0/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1443 comparator_0/xnor_2/not_0/in comparator_0/xnor_2/XOR_0/bbar a1out_2 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1444 comparator_0/a0xnorb0 comparator_0/xnor_3/not_0/in vdd comparator_0/xnor_3/not_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1445 comparator_0/a0xnorb0 comparator_0/xnor_3/not_0/in gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1446 comparator_0/xnor_3/not_0/in boout_2 comparator_0/xnor_3/XOR_0/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1447 comparator_0/xnor_3/XOR_0/bbar boout_2 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1448 comparator_0/xnor_3/not_0/in comparator_0/xnor_3/XOR_0/bbar comparator_0/xnor_3/XOR_0/abar comparator_0/xnor_3/XOR_0/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1449 vdd boout_2 comparator_0/xnor_3/XOR_0/bbar comparator_0/xnor_3/XOR_0/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1450 comparator_0/xnor_3/not_0/in boout_2 a0out_2 comparator_0/xnor_3/XOR_0/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1451 comparator_0/xnor_3/XOR_0/abar a0out_2 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1452 vdd a0out_2 comparator_0/xnor_3/XOR_0/abar comparator_0/xnor_3/XOR_0/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1453 comparator_0/xnor_3/not_0/in comparator_0/xnor_3/XOR_0/bbar a0out_2 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1454 comparator_0/a1bar a1out_2 vdd comparator_0/not_5/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1455 comparator_0/a1bar a1out_2 gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1456 comparator_0/a2bar a2out_2 vdd comparator_0/not_6/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1457 comparator_0/a2bar a2out_2 gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1458 comparator_0/a3bar a3out_2 vdd comparator_0/not_7/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1459 comparator_0/a3bar a3out_2 gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1460 comparator_0/t8 comparator_0/5input_AND_0/not_0/in vdd comparator_0/5input_AND_0/not_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1461 comparator_0/t8 comparator_0/5input_AND_0/not_0/in gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1462 vdd a0out_2 comparator_0/5input_AND_0/not_0/in comparator_0/5input_AND_0/w_n37_15# CMOSP w=14 l=8
+  ad=0 pd=0 as=405 ps=198
M1463 vdd comparator_0/a3xnorb3 comparator_0/5input_AND_0/not_0/in comparator_0/5input_AND_0/w_31_n55# CMOSP w=15 l=8
+  ad=0 pd=0 as=0 ps=0
M1464 comparator_0/5input_AND_0/a_n33_n203# comparator_0/b0bar comparator_0/5input_AND_0/a_n33_n226# Gnd CMOSN w=36 l=12
+  ad=468 pd=98 as=396 ps=94
M1465 comparator_0/5input_AND_0/not_0/in comparator_0/a1xnorb1 comparator_0/5input_AND_0/a_n33_n154# Gnd CMOSN w=36 l=12
+  ad=540 pd=102 as=432 ps=96
M1466 vdd comparator_0/a1xnorb1 comparator_0/5input_AND_0/not_0/in comparator_0/5input_AND_0/w_106_n113# CMOSP w=13 l=8
+  ad=0 pd=0 as=0 ps=0
M1467 comparator_0/5input_AND_0/a_n33_n154# comparator_0/a2xnorb2 comparator_0/5input_AND_0/a_n33_n178# Gnd CMOSN w=36 l=12
+  ad=0 pd=0 as=432 ps=96
M1468 comparator_0/5input_AND_0/a_n33_n178# comparator_0/a3xnorb3 comparator_0/5input_AND_0/a_n33_n203# Gnd CMOSN w=36 l=12
+  ad=0 pd=0 as=0 ps=0
M1469 comparator_0/5input_AND_0/a_n33_n226# a0out_2 gnd Gnd CMOSN w=36 l=12
+  ad=0 pd=0 as=0 ps=0
M1470 vdd comparator_0/b0bar comparator_0/5input_AND_0/not_0/in comparator_0/5input_AND_0/w_n4_n20# CMOSP w=13 l=8
+  ad=0 pd=0 as=0 ps=0
M1471 vdd comparator_0/a2xnorb2 comparator_0/5input_AND_0/not_0/in comparator_0/5input_AND_0/w_68_n82# CMOSP w=14 l=8
+  ad=0 pd=0 as=0 ps=0
M1472 comparator_0/t4 comparator_0/5input_AND_1/not_0/in vdd comparator_0/5input_AND_1/not_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1473 comparator_0/t4 comparator_0/5input_AND_1/not_0/in gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1474 vdd comparator_0/a0bar comparator_0/5input_AND_1/not_0/in comparator_0/5input_AND_1/w_n37_15# CMOSP w=14 l=8
+  ad=0 pd=0 as=405 ps=198
M1475 vdd comparator_0/a1xnorb1 comparator_0/5input_AND_1/not_0/in comparator_0/5input_AND_1/w_31_n55# CMOSP w=15 l=8
+  ad=0 pd=0 as=0 ps=0
M1476 comparator_0/5input_AND_1/a_n33_n203# boout_2 comparator_0/5input_AND_1/a_n33_n226# Gnd CMOSN w=36 l=12
+  ad=468 pd=98 as=396 ps=94
M1477 comparator_0/5input_AND_1/not_0/in comparator_0/a3xnorb3 comparator_0/5input_AND_1/a_n33_n154# Gnd CMOSN w=36 l=12
+  ad=540 pd=102 as=432 ps=96
M1478 vdd comparator_0/a3xnorb3 comparator_0/5input_AND_1/not_0/in comparator_0/5input_AND_1/w_106_n113# CMOSP w=13 l=8
+  ad=0 pd=0 as=0 ps=0
M1479 comparator_0/5input_AND_1/a_n33_n154# comparator_0/a2xnorb2 comparator_0/5input_AND_1/a_n33_n178# Gnd CMOSN w=36 l=12
+  ad=0 pd=0 as=432 ps=96
M1480 comparator_0/5input_AND_1/a_n33_n178# comparator_0/a1xnorb1 comparator_0/5input_AND_1/a_n33_n203# Gnd CMOSN w=36 l=12
+  ad=0 pd=0 as=0 ps=0
M1481 comparator_0/5input_AND_1/a_n33_n226# comparator_0/a0bar gnd Gnd CMOSN w=36 l=12
+  ad=0 pd=0 as=0 ps=0
M1482 vdd boout_2 comparator_0/5input_AND_1/not_0/in comparator_0/5input_AND_1/w_n4_n20# CMOSP w=13 l=8
+  ad=0 pd=0 as=0 ps=0
M1483 vdd comparator_0/a2xnorb2 comparator_0/5input_AND_1/not_0/in comparator_0/5input_AND_1/w_68_n82# CMOSP w=14 l=8
+  ad=0 pd=0 as=0 ps=0
M1484 comparator_0/t5 comparator_0/and_0/a_n26_14# vdd comparator_0/and_0/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1485 vdd comparator_0/b3bar comparator_0/and_0/a_n26_14# comparator_0/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1486 comparator_0/t5 comparator_0/and_0/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1487 comparator_0/and_0/a_n26_14# a3out_2 vdd comparator_0/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1488 comparator_0/and_0/a_n26_n23# a3out_2 gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1489 comparator_0/and_0/a_n26_14# comparator_0/b3bar comparator_0/and_0/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1490 equal comparator_0/4input_AND_0/not_0/in vdd comparator_0/4input_AND_0/not_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1491 equal comparator_0/4input_AND_0/not_0/in gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1492 vdd comparator_0/a3xnorb3 comparator_0/4input_AND_0/not_0/in comparator_0/4input_AND_0/w_n47_52# CMOSP w=12 l=7
+  ad=0 pd=0 as=648 ps=204
M1493 comparator_0/4input_AND_0/not_0/in comparator_0/a0xnorb0 comparator_0/4input_AND_0/a_n40_n132# Gnd CMOSN w=12 l=7
+  ad=120 pd=44 as=96 ps=40
M1494 comparator_0/4input_AND_0/a_n40_n147# comparator_0/a2xnorb2 comparator_0/4input_AND_0/a_n40_n162# Gnd CMOSN w=12 l=7
+  ad=96 pd=40 as=96 ps=40
M1495 vdd comparator_0/a0xnorb0 comparator_0/4input_AND_0/not_0/in comparator_0/4input_AND_0/w_68_n95# CMOSP w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1496 comparator_0/4input_AND_0/a_n40_n132# comparator_0/a1xnorb1 comparator_0/4input_AND_0/a_n40_n147# Gnd CMOSN w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1497 comparator_0/4input_AND_0/a_n40_n162# comparator_0/a3xnorb3 gnd Gnd CMOSN w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1498 vdd comparator_0/a2xnorb2 comparator_0/4input_AND_0/not_0/in comparator_0/4input_AND_0/w_n8_2# CMOSP w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1499 vdd comparator_0/a1xnorb1 comparator_0/4input_AND_0/not_0/in comparator_0/4input_AND_0/w_29_n46# CMOSP w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1500 comparator_0/t7 comparator_0/4input_AND_1/not_0/in vdd comparator_0/4input_AND_1/not_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1501 comparator_0/t7 comparator_0/4input_AND_1/not_0/in gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1502 vdd a1out_2 comparator_0/4input_AND_1/not_0/in comparator_0/4input_AND_1/w_n47_52# CMOSP w=12 l=7
+  ad=0 pd=0 as=648 ps=204
M1503 comparator_0/4input_AND_1/not_0/in comparator_0/a2xnorb2 comparator_0/4input_AND_1/a_n40_n132# Gnd CMOSN w=12 l=7
+  ad=120 pd=44 as=96 ps=40
M1504 comparator_0/4input_AND_1/a_n40_n147# comparator_0/b1bar comparator_0/4input_AND_1/a_n40_n162# Gnd CMOSN w=12 l=7
+  ad=96 pd=40 as=96 ps=40
M1505 vdd comparator_0/a2xnorb2 comparator_0/4input_AND_1/not_0/in comparator_0/4input_AND_1/w_68_n95# CMOSP w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1506 comparator_0/4input_AND_1/a_n40_n132# comparator_0/a3xnorb3 comparator_0/4input_AND_1/a_n40_n147# Gnd CMOSN w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1507 comparator_0/4input_AND_1/a_n40_n162# a1out_2 gnd Gnd CMOSN w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1508 vdd comparator_0/b1bar comparator_0/4input_AND_1/not_0/in comparator_0/4input_AND_1/w_n8_2# CMOSP w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1509 vdd comparator_0/a3xnorb3 comparator_0/4input_AND_1/not_0/in comparator_0/4input_AND_1/w_29_n46# CMOSP w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1510 comparator_0/t1 comparator_0/and_1/a_n26_14# vdd comparator_0/and_1/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1511 vdd b3out_2 comparator_0/and_1/a_n26_14# comparator_0/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1512 comparator_0/t1 comparator_0/and_1/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1513 comparator_0/and_1/a_n26_14# comparator_0/a3bar vdd comparator_0/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1514 comparator_0/and_1/a_n26_n23# comparator_0/a3bar gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1515 comparator_0/and_1/a_n26_14# b3out_2 comparator_0/and_1/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1516 comparator_0/t3 comparator_0/4input_AND_2/not_0/in vdd comparator_0/4input_AND_2/not_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1517 comparator_0/t3 comparator_0/4input_AND_2/not_0/in gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1518 vdd comparator_0/a1bar comparator_0/4input_AND_2/not_0/in comparator_0/4input_AND_2/w_n47_52# CMOSP w=12 l=7
+  ad=0 pd=0 as=648 ps=204
M1519 comparator_0/4input_AND_2/not_0/in comparator_0/a3xnorb3 comparator_0/4input_AND_2/a_n40_n132# Gnd CMOSN w=12 l=7
+  ad=120 pd=44 as=96 ps=40
M1520 comparator_0/4input_AND_2/a_n40_n147# b1out_2 comparator_0/4input_AND_2/a_n40_n162# Gnd CMOSN w=12 l=7
+  ad=96 pd=40 as=96 ps=40
M1521 vdd comparator_0/a3xnorb3 comparator_0/4input_AND_2/not_0/in comparator_0/4input_AND_2/w_68_n95# CMOSP w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1522 comparator_0/4input_AND_2/a_n40_n132# comparator_0/a2xnorb2 comparator_0/4input_AND_2/a_n40_n147# Gnd CMOSN w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1523 comparator_0/4input_AND_2/a_n40_n162# comparator_0/a1bar gnd Gnd CMOSN w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1524 vdd b1out_2 comparator_0/4input_AND_2/not_0/in comparator_0/4input_AND_2/w_n8_2# CMOSP w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1525 vdd comparator_0/a2xnorb2 comparator_0/4input_AND_2/not_0/in comparator_0/4input_AND_2/w_29_n46# CMOSP w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1526 comparator_0/t6 comparator_0/3input_AND_0/not_0/in vdd comparator_0/3input_AND_0/not_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1527 comparator_0/t6 comparator_0/3input_AND_0/not_0/in gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1528 comparator_0/3input_AND_0/a_n9_n125# comparator_0/b2bar gnd Gnd CMOSN w=15 l=8
+  ad=135 pd=48 as=0 ps=0
M1529 comparator_0/3input_AND_0/not_0/in comparator_0/a3xnorb3 comparator_0/3input_AND_0/a_n9_n108# Gnd CMOSN w=15 l=8
+  ad=165 pd=52 as=165 ps=52
M1530 vdd comparator_0/a3xnorb3 comparator_0/3input_AND_0/not_0/in comparator_0/3input_AND_0/w_69_n71# CMOSP w=13 l=8
+  ad=0 pd=0 as=546 ps=162
M1531 vdd a2out_2 comparator_0/3input_AND_0/not_0/in comparator_0/3input_AND_0/w_32_n21# CMOSP w=13 l=8
+  ad=0 pd=0 as=0 ps=0
M1532 vdd comparator_0/b2bar comparator_0/3input_AND_0/not_0/in comparator_0/3input_AND_0/w_n14_24# CMOSP w=13 l=8
+  ad=0 pd=0 as=0 ps=0
M1533 comparator_0/3input_AND_0/a_n9_n108# a2out_2 comparator_0/3input_AND_0/a_n9_n125# Gnd CMOSN w=15 l=8
+  ad=0 pd=0 as=0 ps=0
M1534 comparator_0/t2 comparator_0/3input_AND_1/not_0/in vdd comparator_0/3input_AND_1/not_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1535 comparator_0/t2 comparator_0/3input_AND_1/not_0/in gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1536 comparator_0/3input_AND_1/a_n9_n125# comparator_0/a2bar gnd Gnd CMOSN w=15 l=8
+  ad=135 pd=48 as=0 ps=0
M1537 comparator_0/3input_AND_1/not_0/in comparator_0/a3xnorb3 comparator_0/3input_AND_1/a_n9_n108# Gnd CMOSN w=15 l=8
+  ad=165 pd=52 as=165 ps=52
M1538 vdd comparator_0/a3xnorb3 comparator_0/3input_AND_1/not_0/in comparator_0/3input_AND_1/w_69_n71# CMOSP w=13 l=8
+  ad=0 pd=0 as=546 ps=162
M1539 vdd b2out_2 comparator_0/3input_AND_1/not_0/in comparator_0/3input_AND_1/w_32_n21# CMOSP w=13 l=8
+  ad=0 pd=0 as=0 ps=0
M1540 vdd comparator_0/a2bar comparator_0/3input_AND_1/not_0/in comparator_0/3input_AND_1/w_n14_24# CMOSP w=13 l=8
+  ad=0 pd=0 as=0 ps=0
M1541 comparator_0/3input_AND_1/a_n9_n108# b2out_2 comparator_0/3input_AND_1/a_n9_n125# Gnd CMOSN w=15 l=8
+  ad=0 pd=0 as=0 ps=0
M1542 4bitadder_1/fulladder_0/or_0/a_n15_32# 4bitadder_1/fulladder_0/or_0/a gnd Gnd CMOSN w=16 l=5
+  ad=304 pd=70 as=0 ps=0
M1543 4bitadder_1/c1 4bitadder_1/fulladder_0/or_0/a_n15_32# vdd 4bitadder_1/fulladder_0/or_0/w_58_101# CMOSP w=16 l=6
+  ad=288 pd=68 as=0 ps=0
M1544 gnd 4bitadder_1/fulladder_0/or_0/b 4bitadder_1/fulladder_0/or_0/a_n15_32# Gnd CMOSN w=16 l=5
+  ad=0 pd=0 as=0 ps=0
M1545 4bitadder_1/fulladder_0/or_0/a_n15_32# 4bitadder_1/fulladder_0/or_0/b 4bitadder_1/fulladder_0/or_0/a_n15_107# 4bitadder_1/fulladder_0/or_0/w_n48_101# CMOSP w=16 l=5
+  ad=448 pd=88 as=304 ps=70
M1546 4bitadder_1/c1 4bitadder_1/fulladder_0/or_0/a_n15_32# gnd Gnd CMOSN w=16 l=6
+  ad=320 pd=72 as=0 ps=0
M1547 4bitadder_1/fulladder_0/or_0/a_n15_107# 4bitadder_1/fulladder_0/or_0/a vdd 4bitadder_1/fulladder_0/or_0/w_n48_101# CMOSP w=16 l=5
+  ad=0 pd=0 as=0 ps=0
M1548 4bitadder_1/fulladder_0/or_0/a 4bitadder_1/fulladder_0/and_0/a_n26_14# vdd 4bitadder_1/fulladder_0/and_0/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1549 vdd s0 4bitadder_1/fulladder_0/and_0/a_n26_14# 4bitadder_1/fulladder_0/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1550 4bitadder_1/fulladder_0/or_0/a 4bitadder_1/fulladder_0/and_0/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1551 4bitadder_1/fulladder_0/and_0/a_n26_14# 4bitadder_1/fulladder_0/axorb vdd 4bitadder_1/fulladder_0/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1552 4bitadder_1/fulladder_0/and_0/a_n26_n23# 4bitadder_1/fulladder_0/axorb gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1553 4bitadder_1/fulladder_0/and_0/a_n26_14# s0 4bitadder_1/fulladder_0/and_0/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1554 4bitadder_1/fulladder_0/axorb 4bitadder_1/b0xorM 4bitadder_1/fulladder_0/XOR_0/abar Gnd CMOSN w=11 l=6
+  ad=495 pd=156 as=407 ps=118
M1555 4bitadder_1/fulladder_0/XOR_0/bbar 4bitadder_1/b0xorM gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1556 4bitadder_1/fulladder_0/axorb 4bitadder_1/fulladder_0/XOR_0/bbar 4bitadder_1/fulladder_0/XOR_0/abar 4bitadder_1/fulladder_0/XOR_0/w_62_n20# CMOSP w=12 l=6
+  ad=252 pd=110 as=218 ps=84
M1557 vdd 4bitadder_1/b0xorM 4bitadder_1/fulladder_0/XOR_0/bbar 4bitadder_1/fulladder_0/XOR_0/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1558 4bitadder_1/fulladder_0/axorb 4bitadder_1/b0xorM a0_out1 4bitadder_1/fulladder_0/XOR_0/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1559 4bitadder_1/fulladder_0/XOR_0/abar a0_out1 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1560 vdd a0_out1 4bitadder_1/fulladder_0/XOR_0/abar 4bitadder_1/fulladder_0/XOR_0/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1561 4bitadder_1/fulladder_0/axorb 4bitadder_1/fulladder_0/XOR_0/bbar a0_out1 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1562 4bitadder_1/fulladder_0/or_0/b 4bitadder_1/fulladder_0/and_1/a_n26_14# vdd 4bitadder_1/fulladder_0/and_1/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1563 vdd a0_out1 4bitadder_1/fulladder_0/and_1/a_n26_14# 4bitadder_1/fulladder_0/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1564 4bitadder_1/fulladder_0/or_0/b 4bitadder_1/fulladder_0/and_1/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1565 4bitadder_1/fulladder_0/and_1/a_n26_14# 4bitadder_1/b0xorM vdd 4bitadder_1/fulladder_0/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1566 4bitadder_1/fulladder_0/and_1/a_n26_n23# 4bitadder_1/b0xorM gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1567 4bitadder_1/fulladder_0/and_1/a_n26_14# a0_out1 4bitadder_1/fulladder_0/and_1/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1568 s0_sub s0 4bitadder_1/fulladder_0/XOR_1/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1569 4bitadder_1/fulladder_0/XOR_1/bbar s0 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1570 s0_sub 4bitadder_1/fulladder_0/XOR_1/bbar 4bitadder_1/fulladder_0/XOR_1/abar 4bitadder_1/fulladder_0/XOR_1/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1571 vdd s0 4bitadder_1/fulladder_0/XOR_1/bbar 4bitadder_1/fulladder_0/XOR_1/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1572 s0_sub s0 4bitadder_1/fulladder_0/axorb 4bitadder_1/fulladder_0/XOR_1/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1573 4bitadder_1/fulladder_0/XOR_1/abar 4bitadder_1/fulladder_0/axorb gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1574 vdd 4bitadder_1/fulladder_0/axorb 4bitadder_1/fulladder_0/XOR_1/abar 4bitadder_1/fulladder_0/XOR_1/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1575 s0_sub 4bitadder_1/fulladder_0/XOR_1/bbar 4bitadder_1/fulladder_0/axorb Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1576 4bitadder_1/fulladder_1/or_0/a_n15_32# 4bitadder_1/fulladder_1/or_0/a gnd Gnd CMOSN w=16 l=5
+  ad=304 pd=70 as=0 ps=0
M1577 4bitadder_1/c2 4bitadder_1/fulladder_1/or_0/a_n15_32# vdd 4bitadder_1/fulladder_1/or_0/w_58_101# CMOSP w=16 l=6
+  ad=288 pd=68 as=0 ps=0
M1578 gnd 4bitadder_1/fulladder_1/or_0/b 4bitadder_1/fulladder_1/or_0/a_n15_32# Gnd CMOSN w=16 l=5
+  ad=0 pd=0 as=0 ps=0
M1579 4bitadder_1/fulladder_1/or_0/a_n15_32# 4bitadder_1/fulladder_1/or_0/b 4bitadder_1/fulladder_1/or_0/a_n15_107# 4bitadder_1/fulladder_1/or_0/w_n48_101# CMOSP w=16 l=5
+  ad=448 pd=88 as=304 ps=70
M1580 4bitadder_1/c2 4bitadder_1/fulladder_1/or_0/a_n15_32# gnd Gnd CMOSN w=16 l=6
+  ad=320 pd=72 as=0 ps=0
M1581 4bitadder_1/fulladder_1/or_0/a_n15_107# 4bitadder_1/fulladder_1/or_0/a vdd 4bitadder_1/fulladder_1/or_0/w_n48_101# CMOSP w=16 l=5
+  ad=0 pd=0 as=0 ps=0
M1582 4bitadder_1/fulladder_1/or_0/a 4bitadder_1/fulladder_1/and_0/a_n26_14# vdd 4bitadder_1/fulladder_1/and_0/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1583 vdd 4bitadder_1/c1 4bitadder_1/fulladder_1/and_0/a_n26_14# 4bitadder_1/fulladder_1/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1584 4bitadder_1/fulladder_1/or_0/a 4bitadder_1/fulladder_1/and_0/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1585 4bitadder_1/fulladder_1/and_0/a_n26_14# 4bitadder_1/fulladder_1/axorb vdd 4bitadder_1/fulladder_1/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1586 4bitadder_1/fulladder_1/and_0/a_n26_n23# 4bitadder_1/fulladder_1/axorb gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1587 4bitadder_1/fulladder_1/and_0/a_n26_14# 4bitadder_1/c1 4bitadder_1/fulladder_1/and_0/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1588 4bitadder_1/fulladder_1/axorb 4bitadder_1/XOR_1/out 4bitadder_1/fulladder_1/XOR_0/abar Gnd CMOSN w=11 l=6
+  ad=495 pd=156 as=407 ps=118
M1589 4bitadder_1/fulladder_1/XOR_0/bbar 4bitadder_1/XOR_1/out gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1590 4bitadder_1/fulladder_1/axorb 4bitadder_1/fulladder_1/XOR_0/bbar 4bitadder_1/fulladder_1/XOR_0/abar 4bitadder_1/fulladder_1/XOR_0/w_62_n20# CMOSP w=12 l=6
+  ad=252 pd=110 as=218 ps=84
M1591 vdd 4bitadder_1/XOR_1/out 4bitadder_1/fulladder_1/XOR_0/bbar 4bitadder_1/fulladder_1/XOR_0/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1592 4bitadder_1/fulladder_1/axorb 4bitadder_1/XOR_1/out a1out_1 4bitadder_1/fulladder_1/XOR_0/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1593 4bitadder_1/fulladder_1/XOR_0/abar a1out_1 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1594 vdd a1out_1 4bitadder_1/fulladder_1/XOR_0/abar 4bitadder_1/fulladder_1/XOR_0/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1595 4bitadder_1/fulladder_1/axorb 4bitadder_1/fulladder_1/XOR_0/bbar a1out_1 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1596 4bitadder_1/fulladder_1/or_0/b 4bitadder_1/fulladder_1/and_1/a_n26_14# vdd 4bitadder_1/fulladder_1/and_1/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1597 vdd a1out_1 4bitadder_1/fulladder_1/and_1/a_n26_14# 4bitadder_1/fulladder_1/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1598 4bitadder_1/fulladder_1/or_0/b 4bitadder_1/fulladder_1/and_1/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1599 4bitadder_1/fulladder_1/and_1/a_n26_14# 4bitadder_1/XOR_1/out vdd 4bitadder_1/fulladder_1/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1600 4bitadder_1/fulladder_1/and_1/a_n26_n23# 4bitadder_1/XOR_1/out gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1601 4bitadder_1/fulladder_1/and_1/a_n26_14# a1out_1 4bitadder_1/fulladder_1/and_1/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1602 s1_sub 4bitadder_1/c1 4bitadder_1/fulladder_1/XOR_1/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1603 4bitadder_1/fulladder_1/XOR_1/bbar 4bitadder_1/c1 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1604 s1_sub 4bitadder_1/fulladder_1/XOR_1/bbar 4bitadder_1/fulladder_1/XOR_1/abar 4bitadder_1/fulladder_1/XOR_1/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1605 vdd 4bitadder_1/c1 4bitadder_1/fulladder_1/XOR_1/bbar 4bitadder_1/fulladder_1/XOR_1/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1606 s1_sub 4bitadder_1/c1 4bitadder_1/fulladder_1/axorb 4bitadder_1/fulladder_1/XOR_1/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1607 4bitadder_1/fulladder_1/XOR_1/abar 4bitadder_1/fulladder_1/axorb gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1608 vdd 4bitadder_1/fulladder_1/axorb 4bitadder_1/fulladder_1/XOR_1/abar 4bitadder_1/fulladder_1/XOR_1/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1609 s1_sub 4bitadder_1/fulladder_1/XOR_1/bbar 4bitadder_1/fulladder_1/axorb Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1610 4bitadder_1/fulladder_2/or_0/a_n15_32# 4bitadder_1/fulladder_2/or_0/a gnd Gnd CMOSN w=16 l=5
+  ad=304 pd=70 as=0 ps=0
M1611 4bitadder_1/c3 4bitadder_1/fulladder_2/or_0/a_n15_32# vdd 4bitadder_1/fulladder_2/or_0/w_58_101# CMOSP w=16 l=6
+  ad=288 pd=68 as=0 ps=0
M1612 gnd 4bitadder_1/fulladder_2/or_0/b 4bitadder_1/fulladder_2/or_0/a_n15_32# Gnd CMOSN w=16 l=5
+  ad=0 pd=0 as=0 ps=0
M1613 4bitadder_1/fulladder_2/or_0/a_n15_32# 4bitadder_1/fulladder_2/or_0/b 4bitadder_1/fulladder_2/or_0/a_n15_107# 4bitadder_1/fulladder_2/or_0/w_n48_101# CMOSP w=16 l=5
+  ad=448 pd=88 as=304 ps=70
M1614 4bitadder_1/c3 4bitadder_1/fulladder_2/or_0/a_n15_32# gnd Gnd CMOSN w=16 l=6
+  ad=320 pd=72 as=0 ps=0
M1615 4bitadder_1/fulladder_2/or_0/a_n15_107# 4bitadder_1/fulladder_2/or_0/a vdd 4bitadder_1/fulladder_2/or_0/w_n48_101# CMOSP w=16 l=5
+  ad=0 pd=0 as=0 ps=0
M1616 4bitadder_1/fulladder_2/or_0/a 4bitadder_1/fulladder_2/and_0/a_n26_14# vdd 4bitadder_1/fulladder_2/and_0/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1617 vdd 4bitadder_1/c2 4bitadder_1/fulladder_2/and_0/a_n26_14# 4bitadder_1/fulladder_2/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1618 4bitadder_1/fulladder_2/or_0/a 4bitadder_1/fulladder_2/and_0/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1619 4bitadder_1/fulladder_2/and_0/a_n26_14# 4bitadder_1/fulladder_2/axorb vdd 4bitadder_1/fulladder_2/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1620 4bitadder_1/fulladder_2/and_0/a_n26_n23# 4bitadder_1/fulladder_2/axorb gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1621 4bitadder_1/fulladder_2/and_0/a_n26_14# 4bitadder_1/c2 4bitadder_1/fulladder_2/and_0/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1622 4bitadder_1/fulladder_2/axorb 4bitadder_1/XOR_2/out 4bitadder_1/fulladder_2/XOR_0/abar Gnd CMOSN w=11 l=6
+  ad=495 pd=156 as=407 ps=118
M1623 4bitadder_1/fulladder_2/XOR_0/bbar 4bitadder_1/XOR_2/out gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1624 4bitadder_1/fulladder_2/axorb 4bitadder_1/fulladder_2/XOR_0/bbar 4bitadder_1/fulladder_2/XOR_0/abar 4bitadder_1/fulladder_2/XOR_0/w_62_n20# CMOSP w=12 l=6
+  ad=252 pd=110 as=218 ps=84
M1625 vdd 4bitadder_1/XOR_2/out 4bitadder_1/fulladder_2/XOR_0/bbar 4bitadder_1/fulladder_2/XOR_0/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1626 4bitadder_1/fulladder_2/axorb 4bitadder_1/XOR_2/out a2out_1 4bitadder_1/fulladder_2/XOR_0/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1627 4bitadder_1/fulladder_2/XOR_0/abar a2out_1 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1628 vdd a2out_1 4bitadder_1/fulladder_2/XOR_0/abar 4bitadder_1/fulladder_2/XOR_0/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1629 4bitadder_1/fulladder_2/axorb 4bitadder_1/fulladder_2/XOR_0/bbar a2out_1 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1630 4bitadder_1/fulladder_2/or_0/b 4bitadder_1/fulladder_2/and_1/a_n26_14# vdd 4bitadder_1/fulladder_2/and_1/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1631 vdd a2out_1 4bitadder_1/fulladder_2/and_1/a_n26_14# 4bitadder_1/fulladder_2/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1632 4bitadder_1/fulladder_2/or_0/b 4bitadder_1/fulladder_2/and_1/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1633 4bitadder_1/fulladder_2/and_1/a_n26_14# 4bitadder_1/XOR_2/out vdd 4bitadder_1/fulladder_2/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1634 4bitadder_1/fulladder_2/and_1/a_n26_n23# 4bitadder_1/XOR_2/out gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1635 4bitadder_1/fulladder_2/and_1/a_n26_14# a2out_1 4bitadder_1/fulladder_2/and_1/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1636 s2_sub 4bitadder_1/c2 4bitadder_1/fulladder_2/XOR_1/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1637 4bitadder_1/fulladder_2/XOR_1/bbar 4bitadder_1/c2 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1638 s2_sub 4bitadder_1/fulladder_2/XOR_1/bbar 4bitadder_1/fulladder_2/XOR_1/abar 4bitadder_1/fulladder_2/XOR_1/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1639 vdd 4bitadder_1/c2 4bitadder_1/fulladder_2/XOR_1/bbar 4bitadder_1/fulladder_2/XOR_1/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1640 s2_sub 4bitadder_1/c2 4bitadder_1/fulladder_2/axorb 4bitadder_1/fulladder_2/XOR_1/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1641 4bitadder_1/fulladder_2/XOR_1/abar 4bitadder_1/fulladder_2/axorb gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1642 vdd 4bitadder_1/fulladder_2/axorb 4bitadder_1/fulladder_2/XOR_1/abar 4bitadder_1/fulladder_2/XOR_1/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1643 s2_sub 4bitadder_1/fulladder_2/XOR_1/bbar 4bitadder_1/fulladder_2/axorb Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1644 4bitadder_1/fulladder_3/or_0/a_n15_32# 4bitadder_1/fulladder_3/or_0/a gnd Gnd CMOSN w=16 l=5
+  ad=304 pd=70 as=0 ps=0
M1645 fc_sub 4bitadder_1/fulladder_3/or_0/a_n15_32# vdd 4bitadder_1/fulladder_3/or_0/w_58_101# CMOSP w=16 l=6
+  ad=288 pd=68 as=0 ps=0
M1646 gnd 4bitadder_1/fulladder_3/or_0/b 4bitadder_1/fulladder_3/or_0/a_n15_32# Gnd CMOSN w=16 l=5
+  ad=0 pd=0 as=0 ps=0
M1647 4bitadder_1/fulladder_3/or_0/a_n15_32# 4bitadder_1/fulladder_3/or_0/b 4bitadder_1/fulladder_3/or_0/a_n15_107# 4bitadder_1/fulladder_3/or_0/w_n48_101# CMOSP w=16 l=5
+  ad=448 pd=88 as=304 ps=70
M1648 fc_sub 4bitadder_1/fulladder_3/or_0/a_n15_32# gnd Gnd CMOSN w=16 l=6
+  ad=320 pd=72 as=0 ps=0
M1649 4bitadder_1/fulladder_3/or_0/a_n15_107# 4bitadder_1/fulladder_3/or_0/a vdd 4bitadder_1/fulladder_3/or_0/w_n48_101# CMOSP w=16 l=5
+  ad=0 pd=0 as=0 ps=0
M1650 4bitadder_1/fulladder_3/or_0/a 4bitadder_1/fulladder_3/and_0/a_n26_14# vdd 4bitadder_1/fulladder_3/and_0/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1651 vdd 4bitadder_1/c3 4bitadder_1/fulladder_3/and_0/a_n26_14# 4bitadder_1/fulladder_3/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1652 4bitadder_1/fulladder_3/or_0/a 4bitadder_1/fulladder_3/and_0/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1653 4bitadder_1/fulladder_3/and_0/a_n26_14# 4bitadder_1/fulladder_3/axorb vdd 4bitadder_1/fulladder_3/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1654 4bitadder_1/fulladder_3/and_0/a_n26_n23# 4bitadder_1/fulladder_3/axorb gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1655 4bitadder_1/fulladder_3/and_0/a_n26_14# 4bitadder_1/c3 4bitadder_1/fulladder_3/and_0/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1656 4bitadder_1/fulladder_3/axorb 4bitadder_1/XOR_3/out 4bitadder_1/fulladder_3/XOR_0/abar Gnd CMOSN w=11 l=6
+  ad=495 pd=156 as=407 ps=118
M1657 4bitadder_1/fulladder_3/XOR_0/bbar 4bitadder_1/XOR_3/out gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1658 4bitadder_1/fulladder_3/axorb 4bitadder_1/fulladder_3/XOR_0/bbar 4bitadder_1/fulladder_3/XOR_0/abar 4bitadder_1/fulladder_3/XOR_0/w_62_n20# CMOSP w=12 l=6
+  ad=252 pd=110 as=218 ps=84
M1659 vdd 4bitadder_1/XOR_3/out 4bitadder_1/fulladder_3/XOR_0/bbar 4bitadder_1/fulladder_3/XOR_0/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1660 4bitadder_1/fulladder_3/axorb 4bitadder_1/XOR_3/out a3out_1 4bitadder_1/fulladder_3/XOR_0/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1661 4bitadder_1/fulladder_3/XOR_0/abar a3out_1 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1662 vdd a3out_1 4bitadder_1/fulladder_3/XOR_0/abar 4bitadder_1/fulladder_3/XOR_0/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1663 4bitadder_1/fulladder_3/axorb 4bitadder_1/fulladder_3/XOR_0/bbar a3out_1 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1664 4bitadder_1/fulladder_3/or_0/b 4bitadder_1/fulladder_3/and_1/a_n26_14# vdd 4bitadder_1/fulladder_3/and_1/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1665 vdd a3out_1 4bitadder_1/fulladder_3/and_1/a_n26_14# 4bitadder_1/fulladder_3/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1666 4bitadder_1/fulladder_3/or_0/b 4bitadder_1/fulladder_3/and_1/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1667 4bitadder_1/fulladder_3/and_1/a_n26_14# 4bitadder_1/XOR_3/out vdd 4bitadder_1/fulladder_3/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1668 4bitadder_1/fulladder_3/and_1/a_n26_n23# 4bitadder_1/XOR_3/out gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1669 4bitadder_1/fulladder_3/and_1/a_n26_14# a3out_1 4bitadder_1/fulladder_3/and_1/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1670 s3_sub 4bitadder_1/c3 4bitadder_1/fulladder_3/XOR_1/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1671 4bitadder_1/fulladder_3/XOR_1/bbar 4bitadder_1/c3 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1672 s3_sub 4bitadder_1/fulladder_3/XOR_1/bbar 4bitadder_1/fulladder_3/XOR_1/abar 4bitadder_1/fulladder_3/XOR_1/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1673 vdd 4bitadder_1/c3 4bitadder_1/fulladder_3/XOR_1/bbar 4bitadder_1/fulladder_3/XOR_1/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1674 s3_sub 4bitadder_1/c3 4bitadder_1/fulladder_3/axorb 4bitadder_1/fulladder_3/XOR_1/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1675 4bitadder_1/fulladder_3/XOR_1/abar 4bitadder_1/fulladder_3/axorb gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1676 vdd 4bitadder_1/fulladder_3/axorb 4bitadder_1/fulladder_3/XOR_1/abar 4bitadder_1/fulladder_3/XOR_1/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1677 s3_sub 4bitadder_1/fulladder_3/XOR_1/bbar 4bitadder_1/fulladder_3/axorb Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1678 4bitadder_1/b0xorM s0 4bitadder_1/XOR_0/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1679 4bitadder_1/XOR_0/bbar s0 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1680 4bitadder_1/b0xorM 4bitadder_1/XOR_0/bbar 4bitadder_1/XOR_0/abar 4bitadder_1/XOR_0/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1681 vdd s0 4bitadder_1/XOR_0/bbar 4bitadder_1/XOR_0/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1682 4bitadder_1/b0xorM s0 b0out_1 4bitadder_1/XOR_0/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1683 4bitadder_1/XOR_0/abar b0out_1 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1684 vdd b0out_1 4bitadder_1/XOR_0/abar 4bitadder_1/XOR_0/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1685 4bitadder_1/b0xorM 4bitadder_1/XOR_0/bbar b0out_1 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1686 4bitadder_1/XOR_1/out s0 4bitadder_1/XOR_1/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1687 4bitadder_1/XOR_1/bbar s0 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1688 4bitadder_1/XOR_1/out 4bitadder_1/XOR_1/bbar 4bitadder_1/XOR_1/abar 4bitadder_1/XOR_1/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1689 vdd s0 4bitadder_1/XOR_1/bbar 4bitadder_1/XOR_1/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1690 4bitadder_1/XOR_1/out s0 b1out_1 4bitadder_1/XOR_1/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1691 4bitadder_1/XOR_1/abar b1out_1 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1692 vdd b1out_1 4bitadder_1/XOR_1/abar 4bitadder_1/XOR_1/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1693 4bitadder_1/XOR_1/out 4bitadder_1/XOR_1/bbar b1out_1 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1694 4bitadder_1/XOR_2/out s0 4bitadder_1/XOR_2/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1695 4bitadder_1/XOR_2/bbar s0 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1696 4bitadder_1/XOR_2/out 4bitadder_1/XOR_2/bbar 4bitadder_1/XOR_2/abar 4bitadder_1/XOR_2/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1697 vdd s0 4bitadder_1/XOR_2/bbar 4bitadder_1/XOR_2/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1698 4bitadder_1/XOR_2/out s0 b2out_1 4bitadder_1/XOR_2/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1699 4bitadder_1/XOR_2/abar b2out_1 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1700 vdd b2out_1 4bitadder_1/XOR_2/abar 4bitadder_1/XOR_2/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1701 4bitadder_1/XOR_2/out 4bitadder_1/XOR_2/bbar b2out_1 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1702 4bitadder_1/XOR_3/out s0 4bitadder_1/XOR_3/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1703 4bitadder_1/XOR_3/bbar s0 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1704 4bitadder_1/XOR_3/out 4bitadder_1/XOR_3/bbar 4bitadder_1/XOR_3/abar 4bitadder_1/XOR_3/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1705 vdd s0 4bitadder_1/XOR_3/bbar 4bitadder_1/XOR_3/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1706 4bitadder_1/XOR_3/out s0 b3out_1 4bitadder_1/XOR_3/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=0 ps=0
M1707 4bitadder_1/XOR_3/abar b3out_1 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1708 vdd b3out_1 4bitadder_1/XOR_3/abar 4bitadder_1/XOR_3/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1709 4bitadder_1/XOR_3/out 4bitadder_1/XOR_3/bbar b3out_1 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=0 ps=0
M1710 decoder_0/and_2/a s0 vdd decoder_0/not_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1711 decoder_0/and_2/a s0 gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1712 decoder_0/and_1/b s1 vdd decoder_0/not_1/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1713 decoder_0/and_1/b s1 gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1714 enable_0/en decoder_0/and_0/a_n26_14# vdd decoder_0/and_0/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1715 vdd decoder_0/and_1/b decoder_0/and_0/a_n26_14# decoder_0/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1716 enable_0/en decoder_0/and_0/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1717 decoder_0/and_0/a_n26_14# decoder_0/and_2/a vdd decoder_0/and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1718 decoder_0/and_0/a_n26_n23# decoder_0/and_2/a gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1719 decoder_0/and_0/a_n26_14# decoder_0/and_1/b decoder_0/and_0/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1720 enable_1/en decoder_0/and_1/a_n26_14# vdd decoder_0/and_1/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1721 vdd decoder_0/and_1/b decoder_0/and_1/a_n26_14# decoder_0/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1722 enable_1/en decoder_0/and_1/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1723 decoder_0/and_1/a_n26_14# s0 vdd decoder_0/and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1724 decoder_0/and_1/a_n26_n23# s0 gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1725 decoder_0/and_1/a_n26_14# decoder_0/and_1/b decoder_0/and_1/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1726 enable_2/en decoder_0/and_2/a_n26_14# vdd decoder_0/and_2/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1727 vdd s1 decoder_0/and_2/a_n26_14# decoder_0/and_2/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1728 enable_2/en decoder_0/and_2/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1729 decoder_0/and_2/a_n26_14# decoder_0/and_2/a vdd decoder_0/and_2/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1730 decoder_0/and_2/a_n26_n23# decoder_0/and_2/a gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1731 decoder_0/and_2/a_n26_14# s1 decoder_0/and_2/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1732 enable_3/en decoder_0/and_3/a_n26_14# vdd decoder_0/and_3/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1733 vdd s1 decoder_0/and_3/a_n26_14# decoder_0/and_3/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1734 enable_3/en decoder_0/and_3/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1735 decoder_0/and_3/a_n26_14# s0 vdd decoder_0/and_3/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1736 decoder_0/and_3/a_n26_n23# s0 gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1737 decoder_0/and_3/a_n26_14# s1 decoder_0/and_3/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
C0 4bitadder_1/fulladder_2/XOR_0/w_n34_n1# a2out_1 0.11fF
C1 4bitadder_1/fulladder_2/XOR_0/w_16_n1# 4bitadder_1/XOR_2/out 0.11fF
C2 vdd comparator_0/3input_AND_0/w_32_n21# 0.03fF
C3 s0 decoder_0/and_1/b 0.19fF
C4 AND_Block_0/and_1/a_n26_14# AND_Block_0/and_1/w_n43_8# 0.02fF
C5 enable_1/and_3/w_n43_8# vdd 0.07fF
C6 comparator_0/and_0/w_26_9# comparator_0/and_0/a_n26_14# 0.09fF
C7 comparator_0/and_0/w_n43_8# comparator_0/b3bar 0.09fF
C8 4bitadder_1/XOR_1/out 4bitadder_1/XOR_1/w_62_n20# 0.04fF
C9 4bitadder_0/fulladder_3/and_0/a_n26_14# 4bitadder_0/c3 0.10fF
C10 s0 4bitadder_1/XOR_1/bbar 0.02fF
C11 vdd 4bitadder_1/fulladder_1/or_0/w_n48_101# 0.05fF
C12 4bitadder_1/fulladder_1/or_0/w_n48_101# 4bitadder_1/fulladder_1/or_0/b 0.12fF
C13 4bitadder_0/fulladder_3/axorb 4bitadder_0/fulladder_3/XOR_1/abar 0.13fF
C14 4bitadder_1/fulladder_2/XOR_0/abar 4bitadder_1/XOR_2/out 0.25fF
C15 enable_1/and_3/w_n43_8# a3 0.09fF
C16 b1out_3 b0out_3 24.79fF
C17 decoder_0/not_1/w_n2_10# s1 0.09fF
C18 4bitadder_1/c3 4bitadder_1/XOR_3/out 0.41fF
C19 enable_1/and_0/w_26_9# a0_out1 0.03fF
C20 enable_0/and_0/w_26_9# enable_0/and_0/a_n26_14# 0.09fF
C21 gnd 4bitadder_1/XOR_3/abar 0.20fF
C22 4bitadder_0/XOR_1/w_n34_n1# vdd 0.02fF
C23 4bitadder_0/fulladder_1/and_1/w_n43_8# vdd 0.07fF
C24 enable_3/and_5/w_26_9# b1out_3 0.03fF
C25 comparator_0/t5 comparator_0/t7 0.21fF
C26 comparator_0/a1xnorb1 comparator_0/4input_AND_0/w_29_n46# 0.16fF
C27 a0out_2 gnd 0.56fF
C28 4bitadder_0/fulladder_1/XOR_1/w_62_37# s1_add 0.02fF
C29 enable_2/and_2/w_n43_8# enable_2/and_2/a_n26_14# 0.02fF
C30 4bitadder_0/fulladder_0/or_0/a vdd 0.14fF
C31 4bitadder_0/fulladder_0/XOR_0/w_62_n20# 4bitadder_0/fulladder_0/XOR_0/abar 0.02fF
C32 4bitadder_1/fulladder_2/XOR_1/w_62_n20# 4bitadder_1/fulladder_2/XOR_1/bbar 0.13fF
C33 4bitadder_0/c1 gnd 0.77fF
C34 enable_2/en a2 0.31fF
C35 a1 vdd 0.42fF
C36 gnd 4bitadder_1/fulladder_2/axorb 0.09fF
C37 vdd b3out_1 0.13fF
C38 4bitadder_1/fulladder_3/or_0/w_n48_101# 4bitadder_1/fulladder_3/or_0/a_n15_32# 0.05fF
C39 b3out_0 4bitadder_0/XOR_3/w_62_37# 0.02fF
C40 enable_1/and_2/w_n43_8# enable_1/and_2/a_n26_14# 0.02fF
C41 comparator_0/xnor_1/XOR_0/w_16_n1# b2out_2 0.11fF
C42 4bitadder_0/XOR_1/w_62_37# b1out_0 0.02fF
C43 enable_2/and_4/w_n43_8# vdd 0.07fF
C44 a1 a3 0.31fF
C45 a0 b0 0.37fF
C46 4bitadder_1/fulladder_1/or_0/w_58_101# 4bitadder_1/c2 0.02fF
C47 enable_3/and_1/w_26_9# a1out_3 0.03fF
C48 4bitadder_1/fulladder_1/axorb 4bitadder_1/c1 0.54fF
C49 AND_Block_0/and_2/a_n26_14# AND_Block_0/and_2/w_26_9# 0.09fF
C50 vdd s1_sub 0.19fF
C51 vdd boout_2 0.94fF
C52 b2out_0 4bitadder_0/XOR_2/abar 0.13fF
C53 enable_1/and_5/w_26_9# vdd 0.03fF
C54 b3 vdd 0.34fF
C55 b2out_2 comparator_0/xnor_1/XOR_0/abar 0.30fF
C56 b0out_3 gnd 0.22fF
C57 4bitadder_1/c3 4bitadder_1/fulladder_3/and_0/w_n43_8# 0.09fF
C58 4bitadder_0/fulladder_2/XOR_0/w_n34_n1# a2out_0 0.11fF
C59 4bitadder_0/fulladder_2/XOR_0/w_16_n1# 4bitadder_0/XOR_2/out 0.11fF
C60 enable_0/and_6/a_n26_14# b2 0.31fF
C61 4bitadder_1/fulladder_1/or_0/w_n48_101# 4bitadder_1/fulladder_1/or_0/a_n15_32# 0.05fF
C62 enable_1/and_0/a_n26_14# a0 0.31fF
C63 4bitadder_0/fulladder_1/axorb vdd 0.15fF
C64 b3 a3 0.31fF
C65 enable_3/en b0 0.25fF
C66 out0 gnd 0.01fF
C67 4bitadder_0/XOR_0/bbar s0 0.02fF
C68 4bitadder_0/fulladder_2/XOR_0/abar 4bitadder_0/XOR_2/out 0.25fF
C69 a2out_3 AND_Block_0/and_2/w_n43_8# 0.09fF
C70 4bitadder_1/fulladder_0/XOR_1/abar gnd 0.15fF
C71 4bitadder_0/c3 4bitadder_0/XOR_3/out 0.41fF
C72 enable_1/and_0/w_n43_8# vdd 0.07fF
C73 b0out_3 a3out_3 0.14fF
C74 vdd 4bitadder_1/fulladder_0/XOR_0/w_n34_n1# 0.02fF
C75 a0out_2 comparator_0/a2xnorb2 0.38fF
C76 enable_1/and_1/a_n26_14# a1 0.31fF
C77 comparator_0/b0bar a0out_2 0.25fF
C78 comparator_0/xnor_3/XOR_0/w_62_37# boout_2 0.13fF
C79 AND_Block_0/and_2/w_n43_8# vdd 0.07fF
C80 4bitadder_1/XOR_1/w_62_n20# 4bitadder_1/XOR_1/abar 0.02fF
C81 a1out_0 a2out_0 2.80fF
C82 comparator_0/xnor_0/XOR_0/w_62_37# comparator_0/xnor_0/not_0/in 0.02fF
C83 a3out_0 vdd 0.29fF
C84 gnd 4bitadder_1/fulladder_3/XOR_1/abar 0.15fF
C85 agb vdd 0.04fF
C86 4bitadder_0/fulladder_2/XOR_1/w_62_n20# 4bitadder_0/fulladder_2/XOR_1/bbar 0.13fF
C87 a3out_2 comparator_0/a3xnorb3 0.18fF
C88 comparator_0/5input_AND_1/not_0/in comparator_0/a3xnorb3 0.23fF
C89 AND_Block_0/and_0/w_26_9# vdd 0.03fF
C90 decoder_0/and_0/w_n43_8# decoder_0/and_0/a_n26_14# 0.02fF
C91 b3out_2 comparator_0/xnor_0/XOR_0/bbar 0.02fF
C92 4bitadder_0/fulladder_3/or_0/w_n48_101# 4bitadder_0/fulladder_3/or_0/a_n15_32# 0.05fF
C93 4bitadder_0/fulladder_1/XOR_0/w_n34_n1# vdd 0.02fF
C94 comparator_0/4input_AND_1/w_29_n46# comparator_0/a3xnorb3 0.16fF
C95 vdd comparator_0/5input_AND_0/w_n4_n20# 0.05fF
C96 out3 gnd 0.01fF
C97 enable_3/and_0/w_26_9# enable_3/and_0/a_n26_14# 0.09fF
C98 s0 b3out_1 0.19fF
C99 4bitadder_1/XOR_2/w_16_n1# 4bitadder_1/XOR_2/bbar 0.03fF
C100 4bitadder_1/XOR_2/w_n34_n1# 4bitadder_1/XOR_2/abar 0.03fF
C101 4bitadder_0/fulladder_2/XOR_1/w_16_n1# vdd 0.02fF
C102 enable_2/and_6/w_n43_8# enable_2/en 0.09fF
C103 comparator_0/a0bar comparator_0/a3xnorb3 0.29fF
C104 comparator_0/b1bar a1out_2 0.18fF
C105 enable_1/and_4/w_n43_8# b0 0.09fF
C106 comparator_0/4input_AND_2/not_0/in gnd 0.24fF
C107 vdd comparator_0/a2bar 0.45fF
C108 4bitadder_0/fulladder_1/or_0/a_n15_32# 4bitadder_0/fulladder_1/or_0/b 0.19fF
C109 a2out_3 vdd 0.12fF
C110 4bitadder_0/c3 4bitadder_0/fulladder_3/and_0/w_n43_8# 0.09fF
C111 gnd s1 0.34fF
C112 vdd b0out_1 0.13fF
C113 comparator_0/and_0/a_n26_14# gnd 0.00fF
C114 enable_0/and_1/w_26_9# enable_0/and_1/a_n26_14# 0.09fF
C115 AND_Block_0/and_3/w_26_9# vdd 0.03fF
C116 4bitadder_1/fulladder_3/or_0/w_n48_101# 4bitadder_1/fulladder_3/or_0/b 0.12fF
C117 comparator_0/3input_AND_0/not_0/in gnd 0.21fF
C118 b3out_3 AND_Block_0/and_3/a_n26_14# 0.31fF
C119 enable_2/and_3/w_n43_8# enable_2/and_3/a_n26_14# 0.02fF
C120 4bitadder_0/fulladder_3/or_0/w_58_101# vdd 0.05fF
C121 a0out_0 vdd 0.26fF
C122 enable_0/and_5/w_26_9# b1out_0 0.03fF
C123 4bitadder_1/fulladder_1/XOR_0/w_n34_n1# a1out_1 0.11fF
C124 comparator_0/b3bar comparator_0/a3xnorb3 0.14fF
C125 decoder_0/and_2/w_n43_8# s1 0.09fF
C126 b3out_2 b1out_2 0.48fF
C127 a3out_2 comparator_0/a1xnorb1 0.17fF
C128 comparator_0/a1xnorb1 comparator_0/5input_AND_1/not_0/in 0.23fF
C129 vdd 4bitadder_1/fulladder_0/axorb 0.15fF
C130 enable_2/en b0 0.31fF
C131 comparator_0/4input_AND_2/w_68_n95# comparator_0/a3xnorb3 0.16fF
C132 AND_Block_0/and_1/w_n43_8# a1out_3 0.09fF
C133 a3 vdd 0.44fF
C134 enable_1/and_3/w_n43_8# enable_1/and_3/a_n26_14# 0.02fF
C135 4bitadder_1/fulladder_3/XOR_0/w_16_n1# 4bitadder_1/fulladder_3/XOR_0/bbar 0.03fF
C136 4bitadder_1/fulladder_3/XOR_0/w_n34_n1# 4bitadder_1/fulladder_3/XOR_0/abar 0.03fF
C137 enable_2/and_5/w_n43_8# b1 0.09fF
C138 comparator_0/4input_AND_1/w_68_n95# comparator_0/a2xnorb2 0.16fF
C139 4bitadder_0/XOR_1/w_62_n20# 4bitadder_0/XOR_1/abar 0.02fF
C140 vdd 4bitadder_1/fulladder_0/and_1/w_26_9# 0.03fF
C141 comparator_0/a0bar comparator_0/a1xnorb1 0.03fF
C142 4bitadder_0/c1 4bitadder_0/fulladder_1/XOR_1/bbar 0.02fF
C143 a2 b0 0.37fF
C144 comparator_0/3input_AND_1/not_0/in comparator_0/3input_AND_1/not_0/w_n2_10# 0.09fF
C145 vdd bga 0.04fF
C146 a2out_2 comparator_0/not_6/w_n2_10# 0.09fF
C147 comparator_0/xnor_1/not_0/w_n2_10# comparator_0/a2xnorb2 0.03fF
C148 a3out_0 s0 0.08fF
C149 vdd comparator_0/t6 0.04fF
C150 comparator_0/4input_AND_2/not_0/in comparator_0/4input_AND_2/w_n8_2# 0.02fF
C151 4bitadder_0/XOR_1/w_n34_n1# b1out_0 0.11fF
C152 b1out_1 b3out_1 0.25fF
C153 decoder_0/and_3/w_n43_8# decoder_0/and_3/a_n26_14# 0.02fF
C154 a1out_2 b1out_2 0.88fF
C155 comparator_0/xnor_2/XOR_0/w_16_n1# comparator_0/xnor_2/XOR_0/bbar 0.03fF
C156 comparator_0/xnor_2/XOR_0/w_62_n20# comparator_0/xnor_2/not_0/in 0.04fF
C157 comparator_0/xnor_2/XOR_0/w_n34_n1# comparator_0/xnor_2/XOR_0/abar 0.03fF
C158 4bitadder_0/fulladder_0/or_0/w_n48_101# 4bitadder_0/fulladder_0/or_0/a_n15_32# 0.05fF
C159 4bitadder_0/XOR_2/w_16_n1# 4bitadder_0/XOR_2/bbar 0.03fF
C160 4bitadder_0/XOR_2/w_n34_n1# 4bitadder_0/XOR_2/abar 0.03fF
C161 4bitadder_0/fulladder_2/or_0/b gnd 0.37fF
C162 comparator_0/4input_AND_2/not_0/in comparator_0/a2xnorb2 0.18fF
C163 4bitadder_1/fulladder_0/and_0/w_26_9# 4bitadder_1/fulladder_0/or_0/a 0.03fF
C164 enable_1/and_5/w_26_9# b1out_1 0.03fF
C165 a3out_1 b2out_1 0.05fF
C166 4bitadder_1/fulladder_1/XOR_0/bbar 4bitadder_1/fulladder_1/XOR_0/w_62_n20# 0.13fF
C167 b0out_0 4bitadder_0/XOR_0/w_n34_n1# 0.11fF
C168 enable_1/and_2/a_n26_14# a2 0.31fF
C169 b0out_0 a1out_0 0.11fF
C170 a0_out1 4bitadder_1/fulladder_0/and_1/w_n43_8# 0.09fF
C171 4bitadder_0/fulladder_3/or_0/w_n48_101# 4bitadder_0/fulladder_3/or_0/b 0.12fF
C172 4bitadder_0/fulladder_2/and_1/w_26_9# vdd 0.03fF
C173 4bitadder_0/fulladder_1/and_1/w_n43_8# 4bitadder_0/fulladder_1/and_1/a_n26_14# 0.02fF
C174 b0out_1 s0 0.17fF
C175 4bitadder_1/fulladder_1/or_0/a_n15_32# 4bitadder_1/fulladder_1/or_0/b 0.19fF
C176 a2out_1 4bitadder_1/fulladder_2/and_1/a_n26_14# 0.10fF
C177 decoder_0/and_1/a_n26_14# decoder_0/and_1/b 0.29fF
C178 vdd decoder_0/and_1/w_26_9# 0.03fF
C179 comparator_0/a1xnorb1 comparator_0/xnor_2/not_0/w_n2_10# 0.03fF
C180 4bitadder_1/fulladder_3/axorb 4bitadder_1/fulladder_3/XOR_1/w_62_37# 0.02fF
C181 4bitadder_1/c3 4bitadder_1/fulladder_3/XOR_1/w_16_n1# 0.11fF
C182 4bitadder_0/fulladder_2/and_0/a_n26_14# 4bitadder_0/fulladder_2/and_0/w_26_9# 0.09fF
C183 vdd s0 0.73fF
C184 4bitadder_1/fulladder_0/XOR_0/w_62_n20# 4bitadder_1/fulladder_0/axorb 0.04fF
C185 a0out_0 s0 0.55fF
C186 gnd decoder_0/and_2/a 0.18fF
C187 comparator_0/a1bar comparator_0/a2xnorb2 0.26fF
C188 b2out_2 comparator_0/3input_AND_1/w_32_n21# 0.16fF
C189 enable_1/and_0/a_n26_14# enable_1/and_0/w_26_9# 0.09fF
C190 a3out_2 b2out_2 0.30fF
C191 b3out_2 a2out_2 0.48fF
C192 comparator_0/5input_AND_1/not_0/in comparator_0/5input_AND_1/w_n4_n20# 0.03fF
C193 4bitadder_1/fulladder_0/axorb s0 0.54fF
C194 4bitadder_0/fulladder_3/XOR_0/w_16_n1# 4bitadder_0/fulladder_3/XOR_0/bbar 0.03fF
C195 4bitadder_0/fulladder_3/XOR_0/w_n34_n1# 4bitadder_0/fulladder_3/XOR_0/abar 0.03fF
C196 AND_Block_0/and_1/a_n26_14# b1out_3 0.31fF
C197 vdd 4bitadder_1/fulladder_2/XOR_1/w_n34_n1# 0.02fF
C198 enable_3/and_1/w_26_9# enable_3/and_1/a_n26_14# 0.09fF
C199 4bitadder_1/c3 4bitadder_1/fulladder_3/XOR_1/abar 0.27fF
C200 4bitadder_1/XOR_1/out a1out_1 1.87fF
C201 comparator_0/not_2/w_n2_10# vdd 0.18fF
C202 decoder_0/and_2/w_n43_8# decoder_0/and_2/a 0.09fF
C203 4bitadder_1/fulladder_3/and_0/a_n26_14# 4bitadder_1/fulladder_3/and_0/w_n43_8# 0.02fF
C204 b3out_0 gnd 0.70fF
C205 b2out_0 a2out_0 0.30fF
C206 b3out_1 4bitadder_1/XOR_3/abar 0.13fF
C207 4bitadder_1/c2 a2out_1 0.50fF
C208 a3out_0 b1out_0 0.12fF
C209 comparator_0/4input_OR_0/w_n58_n43# vdd 0.03fF
C210 enable_0/and_2/w_26_9# enable_0/and_2/a_n26_14# 0.09fF
C211 enable_2/and_4/w_n43_8# enable_2/and_4/a_n26_14# 0.02fF
C212 vdd 4bitadder_1/fulladder_3/and_0/w_n43_8# 0.07fF
C213 4bitadder_1/b0xorM gnd 0.42fF
C214 enable_0/and_7/w_26_9# vdd 0.03fF
C215 a2out_2 a1out_2 0.75fF
C216 4bitadder_1/fulladder_1/XOR_1/w_62_n20# 4bitadder_1/fulladder_1/XOR_1/abar 0.02fF
C217 a0out_2 boout_2 0.87fF
C218 comparator_0/t8 comparator_0/t7 0.15fF
C219 comparator_0/xnor_3/XOR_0/w_16_n1# comparator_0/xnor_3/XOR_0/bbar 0.03fF
C220 comparator_0/xnor_3/XOR_0/w_62_n20# comparator_0/xnor_3/not_0/in 0.04fF
C221 enable_1/en b1 0.25fF
C222 comparator_0/b2bar gnd 0.14fF
C223 comparator_0/3input_AND_1/not_0/in comparator_0/3input_AND_1/w_n14_24# 0.03fF
C224 b2 enable_3/and_6/a_n26_14# 0.31fF
C225 4bitadder_1/fulladder_3/and_1/w_26_9# 4bitadder_1/fulladder_3/and_1/a_n26_14# 0.09fF
C226 enable_1/and_4/w_n43_8# enable_1/and_4/a_n26_14# 0.02fF
C227 enable_2/and_5/w_26_9# b1out_2 0.03fF
C228 comparator_0/4input_AND_0/w_n47_52# comparator_0/a3xnorb3 0.16fF
C229 comparator_0/4input_OR_0/w_n58_n43# comparator_0/t6 0.13fF
C230 vdd b1out_1 0.13fF
C231 gnd 4bitadder_1/fulladder_3/XOR_0/abar 0.15fF
C232 comparator_0/a1xnorb1 comparator_0/5input_AND_1/w_31_n55# 0.21fF
C233 a2out_0 4bitadder_0/fulladder_2/and_1/a_n26_14# 0.10fF
C234 decoder_0/not_0/w_n2_10# decoder_0/and_2/a 0.03fF
C235 comparator_0/3input_AND_1/not_0/in comparator_0/a3xnorb3 0.19fF
C236 vdd 4bitadder_1/fulladder_1/and_0/w_n43_8# 0.07fF
C237 4bitadder_1/XOR_3/out s0 0.16fF
C238 comparator_0/5input_AND_1/w_68_n82# comparator_0/a2xnorb2 0.16fF
C239 4bitadder_0/fulladder_3/axorb 4bitadder_0/fulladder_3/XOR_1/w_62_37# 0.02fF
C240 4bitadder_0/c3 4bitadder_0/fulladder_3/XOR_1/w_16_n1# 0.11fF
C241 4bitadder_0/c1 4bitadder_0/fulladder_1/axorb 0.54fF
C242 4bitadder_1/fulladder_2/XOR_0/w_62_37# 4bitadder_1/XOR_2/out 0.13fF
C243 vdd 4bitadder_1/fulladder_0/XOR_1/w_16_n1# 0.02fF
C244 enable_0/en enable_0/and_6/w_n43_8# 0.09fF
C245 4bitadder_0/XOR_2/abar gnd 0.13fF
C246 4bitadder_1/XOR_1/out 4bitadder_1/fulladder_1/XOR_0/w_62_37# 0.13fF
C247 4bitadder_0/XOR_0/abar gnd 0.15fF
C248 vdd comparator_0/4input_AND_0/w_68_n95# 0.02fF
C249 4bitadder_0/fulladder_2/XOR_0/w_16_n1# vdd 0.02fF
C250 4bitadder_0/XOR_1/out gnd 0.42fF
C251 decoder_0/and_1/b decoder_0/and_1/w_n43_8# 0.09fF
C252 vdd b1out_0 0.13fF
C253 4bitadder_0/c3 4bitadder_0/fulladder_3/XOR_1/abar 0.27fF
C254 comparator_0/t1 gnd 0.01fF
C255 4bitadder_0/fulladder_3/and_0/a_n26_14# 4bitadder_0/fulladder_3/and_0/w_n43_8# 0.02fF
C256 4bitadder_0/fulladder_1/XOR_0/abar a1out_0 0.13fF
C257 4bitadder_1/b0xorM 4bitadder_1/fulladder_0/XOR_0/w_62_37# 0.13fF
C258 b2 a0 0.31fF
C259 4bitadder_0/c2 a2out_0 0.50fF
C260 4bitadder_0/XOR_1/w_16_n1# vdd 0.02fF
C261 4bitadder_1/fulladder_3/or_0/w_n48_101# 4bitadder_1/fulladder_3/or_0/a 0.12fF
C262 comparator_0/3input_AND_0/not_0/in comparator_0/3input_AND_0/w_32_n21# 0.02fF
C263 enable_1/and_3/a_n26_14# a3 0.31fF
C264 vdd 4bitadder_1/fulladder_2/and_1/w_n43_8# 0.07fF
C265 4bitadder_0/fulladder_0/XOR_0/w_16_n1# 4bitadder_0/fulladder_0/XOR_0/bbar 0.03fF
C266 4bitadder_0/fulladder_0/XOR_0/w_n34_n1# 4bitadder_0/fulladder_0/XOR_0/abar 0.03fF
C267 comparator_0/4input_AND_0/w_n8_2# comparator_0/a2xnorb2 0.16fF
C268 enable_1/and_5/w_n43_8# vdd 0.07fF
C269 decoder_0/and_1/b decoder_0/and_2/a 0.34fF
C270 comparator_0/a2xnorb2 comparator_0/b2bar 0.11fF
C271 gnd 4bitadder_1/c2 0.97fF
C272 4bitadder_1/fulladder_1/axorb 4bitadder_1/fulladder_1/XOR_0/w_62_n20# 0.04fF
C273 comparator_0/a0xnorb0 comparator_0/4input_AND_0/not_0/in 0.18fF
C274 comparator_0/xnor_3/XOR_0/abar gnd 0.14fF
C275 vdd 4bitadder_1/XOR_3/w_16_n1# 0.02fF
C276 4bitadder_0/fulladder_1/XOR_1/w_62_n20# 4bitadder_0/fulladder_1/XOR_1/abar 0.02fF
C277 b2 enable_3/en 0.23fF
C278 4bitadder_1/fulladder_2/axorb 4bitadder_1/fulladder_2/XOR_0/w_62_n20# 0.04fF
C279 b2out_0 4bitadder_0/XOR_2/w_62_37# 0.02fF
C280 comparator_0/xnor_1/XOR_0/w_62_37# b2out_2 0.13fF
C281 4bitadder_0/fulladder_3/and_1/w_26_9# 4bitadder_0/fulladder_3/and_1/a_n26_14# 0.09fF
C282 enable_3/and_2/w_26_9# enable_3/and_2/a_n26_14# 0.09fF
C283 b1 gnd 0.27fF
C284 4bitadder_1/fulladder_0/XOR_0/abar a0_out1 0.13fF
C285 vdd a0out_2 0.68fF
C286 b1out_1 s0 0.18fF
C287 b2out_2 comparator_0/xnor_1/not_0/in 0.13fF
C288 a2out_2 comparator_0/xnor_1/XOR_0/abar 0.13fF
C289 4bitadder_0/fulladder_0/and_0/w_n43_8# 4bitadder_0/fulladder_0/and_0/a_n26_14# 0.02fF
C290 4bitadder_0/fulladder_2/XOR_0/w_62_37# 4bitadder_0/XOR_2/out 0.13fF
C291 a0_out1 4bitadder_1/fulladder_0/and_1/a_n26_14# 0.10fF
C292 comparator_0/4input_OR_1/w_n58_n43# comparator_0/t1 0.13fF
C293 4bitadder_0/c1 vdd 0.12fF
C294 enable_0/and_0/w_n43_8# a0 0.09fF
C295 comparator_0/5input_AND_0/not_0/w_n2_10# comparator_0/t8 0.03fF
C296 out0 AND_Block_0/and_0/w_26_9# 0.03fF
C297 enable_0/and_3/w_26_9# enable_0/and_3/a_n26_14# 0.09fF
C298 vdd 4bitadder_1/fulladder_2/axorb 0.15fF
C299 4bitadder_1/fulladder_0/XOR_1/w_16_n1# s0 0.11fF
C300 4bitadder_0/fulladder_2/or_0/a gnd 0.01fF
C301 4bitadder_0/XOR_1/out 4bitadder_0/XOR_1/w_62_37# 0.02fF
C302 a2out_3 b0out_3 0.16fF
C303 s0 b1out_0 13.84fF
C304 4bitadder_1/fulladder_2/or_0/a_n15_32# 4bitadder_1/fulladder_2/or_0/b 0.19fF
C305 comparator_0/5input_AND_0/not_0/in gnd 0.10fF
C306 AND_Block_0/and_0/w_n43_8# vdd 0.07fF
C307 comparator_0/5input_AND_0/not_0/in comparator_0/5input_AND_0/w_68_n82# 0.02fF
C308 enable_0/and_0/w_26_9# vdd 0.03fF
C309 enable_0/and_0/w_26_9# a0out_0 0.03fF
C310 enable_3/and_6/w_n43_8# vdd 0.07fF
C311 4bitadder_1/fulladder_1/and_1/w_n43_8# 4bitadder_1/fulladder_1/and_1/a_n26_14# 0.02fF
C312 4bitadder_1/fulladder_0/or_0/a_n15_32# 4bitadder_1/fulladder_0/or_0/b 0.19fF
C313 4bitadder_0/fulladder_3/or_0/w_n48_101# 4bitadder_0/fulladder_3/or_0/a 0.12fF
C314 a1out_3 b1out_3 2.06fF
C315 comparator_0/xnor_3/XOR_0/w_62_37# a0out_2 0.02fF
C316 b0out_3 vdd 0.16fF
C317 comparator_0/xnor_0/XOR_0/w_n34_n1# a3out_2 0.11fF
C318 4bitadder_0/XOR_1/w_16_n1# s0 0.11fF
C319 a1out_1 enable_1/and_1/w_26_9# 0.03fF
C320 4bitadder_1/fulladder_2/XOR_0/w_62_n20# 4bitadder_1/fulladder_2/XOR_0/bbar 0.13fF
C321 enable_3/and_5/w_26_9# vdd 0.03fF
C322 4bitadder_1/fulladder_3/axorb 4bitadder_1/fulladder_3/XOR_0/w_62_37# 0.02fF
C323 gnd comparator_0/a3xnorb3 0.82fF
C324 b2out_2 comparator_0/3input_AND_1/not_0/in 0.19fF
C325 comparator_0/xnor_3/not_0/w_n2_10# comparator_0/xnor_3/not_0/in 0.09fF
C326 4bitadder_0/fulladder_0/axorb 4bitadder_0/b0xorM 0.13fF
C327 4bitadder_1/XOR_1/out gnd 0.42fF
C328 comparator_0/4input_OR_0/y comparator_0/t7 0.18fF
C329 enable_0/en enable_0/and_1/w_n43_8# 0.09fF
C330 comparator_0/xnor_0/XOR_0/w_62_n20# comparator_0/xnor_0/XOR_0/abar 0.02fF
C331 4bitadder_0/fulladder_3/axorb gnd 0.09fF
C332 4bitadder_0/fulladder_2/axorb 4bitadder_0/fulladder_2/XOR_0/w_62_n20# 0.04fF
C333 vdd 4bitadder_1/fulladder_2/XOR_0/w_n34_n1# 0.02fF
C334 s0 4bitadder_1/XOR_3/w_16_n1# 0.11fF
C335 enable_3/and_0/w_n43_8# a0 0.09fF
C336 b3out_3 gnd 0.24fF
C337 vdd 4bitadder_1/fulladder_3/XOR_1/w_16_n1# 0.02fF
C338 4bitadder_1/fulladder_0/XOR_1/abar 4bitadder_1/fulladder_0/axorb 0.13fF
C339 enable_2/en b2 0.29fF
C340 decoder_0/and_0/w_n43_8# decoder_0/and_1/b 0.09fF
C341 vdd comparator_0/3input_AND_1/w_69_n71# 0.03fF
C342 4bitadder_0/fulladder_1/and_0/w_26_9# 4bitadder_0/fulladder_1/or_0/a 0.03fF
C343 comparator_0/xnor_0/not_0/w_n2_10# comparator_0/xnor_0/not_0/in 0.09fF
C344 comparator_0/4input_AND_0/not_0/w_n2_10# comparator_0/4input_AND_0/not_0/in 0.09fF
C345 s0 4bitadder_1/XOR_3/abar 0.30fF
C346 gnd 4bitadder_1/fulladder_0/or_0/a 0.01fF
C347 s2_add vdd 0.19fF
C348 enable_3/and_0/w_26_9# vdd 0.03fF
C349 enable_2/and_6/w_n43_8# enable_2/and_6/a_n26_14# 0.02fF
C350 vdd comparator_0/4input_AND_1/w_68_n95# 0.02fF
C351 b2 a2 0.31fF
C352 a1out_3 gnd 0.18fF
C353 enable_3/en enable_3/and_0/w_n43_8# 0.09fF
C354 b0out_1 4bitadder_1/XOR_0/w_n34_n1# 0.11fF
C355 enable_1/and_4/a_n26_14# b0 0.31fF
C356 4bitadder_0/fulladder_0/axorb 4bitadder_0/fulladder_0/and_0/w_n43_8# 0.09fF
C357 vdd comparator_0/xnor_1/not_0/w_n2_10# 0.18fF
C358 a3out_3 b3out_3 0.29fF
C359 AND_Block_0/and_3/w_26_9# out3 0.03fF
C360 comparator_0/t4 comparator_0/t3 0.19fF
C361 comparator_0/4input_AND_0/not_0/in comparator_0/4input_AND_0/w_29_n46# 0.02fF
C362 comparator_0/b0bar comparator_0/5input_AND_0/not_0/in 0.23fF
C363 comparator_0/5input_AND_0/not_0/in comparator_0/a2xnorb2 0.23fF
C364 enable_0/and_5/w_n43_8# enable_0/and_5/a_n26_14# 0.02fF
C365 comparator_0/xnor_0/not_0/w_n2_10# vdd 0.18fF
C366 4bitadder_0/fulladder_0/and_1/w_26_9# 4bitadder_0/fulladder_0/and_1/a_n26_14# 0.09fF
C367 vdd 4bitadder_1/XOR_0/w_n34_n1# 0.02fF
C368 a3out_2 b1out_2 0.60fF
C369 comparator_0/a1xnorb1 gnd 1.03fF
C370 b3out_2 a1out_2 0.82fF
C371 4bitadder_1/fulladder_2/axorb 4bitadder_1/fulladder_2/XOR_1/w_n34_n1# 0.11fF
C372 4bitadder_0/fulladder_2/XOR_0/w_62_n20# 4bitadder_0/fulladder_2/XOR_0/bbar 0.13fF
C373 comparator_0/b0bar comparator_0/a3xnorb3 0.28fF
C374 comparator_0/a2xnorb2 comparator_0/a3xnorb3 7.69fF
C375 enable_3/and_3/w_26_9# enable_3/and_3/a_n26_14# 0.09fF
C376 4bitadder_0/fulladder_3/axorb 4bitadder_0/fulladder_3/XOR_0/w_62_37# 0.02fF
C377 4bitadder_0/fulladder_1/or_0/a_n15_32# 4bitadder_0/fulladder_1/or_0/w_58_101# 0.13fF
C378 enable_0/and_6/w_n43_8# vdd 0.07fF
C379 vdd 4bitadder_1/fulladder_2/or_0/w_n48_101# 0.05fF
C380 comparator_0/4input_OR_1/y comparator_0/t3 0.18fF
C381 enable_0/and_1/w_n43_8# a1 0.09fF
C382 comparator_0/t7 comparator_0/4input_AND_1/not_0/w_n2_10# 0.03fF
C383 comparator_0/xnor_2/XOR_0/w_16_n1# b1out_2 0.11fF
C384 4bitadder_0/b0xorM 4bitadder_0/XOR_0/w_62_n20# 0.04fF
C385 enable_0/and_4/w_26_9# enable_0/and_4/a_n26_14# 0.09fF
C386 a2out_0 gnd 1.02fF
C387 gnd 4bitadder_1/fulladder_3/or_0/b 0.37fF
C388 4bitadder_1/fulladder_0/XOR_1/abar s0 0.27fF
C389 vdd comparator_0/a1bar 0.22fF
C390 b1out_2 comparator_0/xnor_2/XOR_0/abar 0.30fF
C391 enable_0/and_2/w_26_9# vdd 0.03fF
C392 gnd 4bitadder_1/XOR_1/abar 0.23fF
C393 comparator_0/4input_AND_2/w_29_n46# comparator_0/a2xnorb2 0.16fF
C394 enable_0/en b1 0.34fF
C395 4bitadder_0/fulladder_1/and_1/w_n43_8# 4bitadder_0/XOR_1/out 0.09fF
C396 comparator_0/a1xnorb1 comparator_0/a2xnorb2 1.39fF
C397 vdd 4bitadder_1/fulladder_3/and_1/w_26_9# 0.03fF
C398 comparator_0/b0bar comparator_0/a1xnorb1 0.29fF
C399 decoder_0/and_1/a_n26_14# decoder_0/and_1/w_26_9# 0.09fF
C400 4bitadder_1/XOR_2/out a2out_1 1.88fF
C401 4bitadder_1/fulladder_2/and_1/w_26_9# 4bitadder_1/fulladder_2/or_0/b 0.03fF
C402 enable_2/and_6/w_n43_8# b2 0.09fF
C403 4bitadder_1/c3 4bitadder_1/fulladder_3/XOR_1/w_62_37# 0.13fF
C404 gnd 4bitadder_1/fulladder_0/or_0/b 0.37fF
C405 4bitadder_1/fulladder_0/XOR_0/w_62_n20# 4bitadder_1/fulladder_0/XOR_0/bbar 0.13fF
C406 4bitadder_0/fulladder_1/XOR_1/abar gnd 0.15fF
C407 4bitadder_0/XOR_3/w_n34_n1# vdd 0.02fF
C408 b2out_2 gnd 0.98fF
C409 enable_0/en enable_0/and_3/w_n43_8# 0.09fF
C410 4bitadder_0/fulladder_2/axorb 4bitadder_0/fulladder_2/XOR_1/w_n34_n1# 0.11fF
C411 b3out_0 a3out_0 0.11fF
C412 a3out_2 a2out_2 0.63fF
C413 vdd decoder_0/and_1/w_n43_8# 0.07fF
C414 a2out_3 enable_3/and_2/w_26_9# 0.03fF
C415 enable_3/and_1/w_n43_8# a1 0.09fF
C416 4bitadder_1/XOR_3/w_62_37# b3out_1 0.02fF
C417 4bitadder_1/c3 s3_sub 0.04fF
C418 4bitadder_0/fulladder_2/and_0/w_26_9# vdd 0.03fF
C419 s0 s1 1.27fF
C420 vdd comparator_0/xnor_1/XOR_0/w_n34_n1# 0.02fF
C421 enable_3/and_2/w_26_9# vdd 0.03fF
C422 4bitadder_1/c1 a1out_1 0.36fF
C423 4bitadder_1/XOR_3/w_62_n20# 4bitadder_1/XOR_3/bbar 0.13fF
C424 b2 b0 0.34fF
C425 enable_3/en enable_3/and_2/w_n43_8# 0.09fF
C426 4bitadder_1/fulladder_0/XOR_1/bbar s0 0.02fF
C427 4bitadder_0/fulladder_3/or_0/w_n48_101# vdd 0.05fF
C428 4bitadder_0/fulladder_1/axorb 4bitadder_0/XOR_1/out 0.13fF
C429 4bitadder_1/fulladder_1/and_1/w_26_9# 4bitadder_1/fulladder_1/and_1/a_n26_14# 0.09fF
C430 vdd decoder_0/and_2/a 0.04fF
C431 vdd comparator_0/5input_AND_1/w_68_n82# 0.05fF
C432 a3out_2 comparator_0/not_7/w_n2_10# 0.09fF
C433 a2out_2 comparator_0/b3bar 0.21fF
C434 4bitadder_1/fulladder_1/XOR_1/w_16_n1# 4bitadder_1/fulladder_1/XOR_1/bbar 0.03fF
C435 4bitadder_1/fulladder_1/XOR_1/w_62_n20# s1_sub 0.04fF
C436 4bitadder_1/fulladder_1/XOR_1/w_n34_n1# 4bitadder_1/fulladder_1/XOR_1/abar 0.03fF
C437 comparator_0/xnor_3/XOR_0/w_16_n1# boout_2 0.11fF
C438 vdd 4bitadder_1/fulladder_1/XOR_0/w_16_n1# 0.02fF
C439 a0_out1 a1out_1 1.88fF
C440 4bitadder_0/fulladder_0/and_0/w_26_9# 4bitadder_0/fulladder_0/or_0/a 0.03fF
C441 4bitadder_1/fulladder_3/and_1/w_n43_8# a3out_1 0.09fF
C442 b3out_0 vdd 0.13fF
C443 b1 a1 0.28fF
C444 decoder_0/and_2/a_n26_14# s1 0.31fF
C445 boout_2 comparator_0/xnor_3/XOR_0/abar 0.30fF
C446 4bitadder_0/XOR_2/out a2out_0 1.88fF
C447 4bitadder_0/fulladder_2/and_1/w_26_9# 4bitadder_0/fulladder_2/or_0/b 0.03fF
C448 enable_3/and_4/w_26_9# enable_3/and_4/a_n26_14# 0.09fF
C449 enable_1/en enable_1/and_2/w_n43_8# 0.09fF
C450 vdd comparator_0/and_0/w_n43_8# 0.07fF
C451 comparator_0/t4 comparator_0/t2 0.19fF
C452 comparator_0/4input_AND_1/not_0/in comparator_0/4input_AND_1/w_29_n46# 0.02fF
C453 enable_0/and_1/w_n43_8# vdd 0.07fF
C454 4bitadder_0/c3 4bitadder_0/fulladder_3/XOR_1/w_62_37# 0.13fF
C455 b0out_0 gnd 0.15fF
C456 4bitadder_0/fulladder_1/XOR_0/w_62_37# a1out_0 0.02fF
C457 b3 b1 0.37fF
C458 4bitadder_1/b0xorM 4bitadder_1/fulladder_0/axorb 0.13fF
C459 vdd comparator_0/4input_AND_0/w_n8_2# 0.02fF
C460 enable_0/and_2/w_n43_8# a2 0.09fF
C461 vdd 4bitadder_1/fulladder_3/XOR_0/w_16_n1# 0.02fF
C462 gnd 4bitadder_1/XOR_2/out 0.42fF
C463 4bitadder_0/c3 s3_add 0.04fF
C464 4bitadder_0/fulladder_1/axorb 4bitadder_0/fulladder_1/and_0/w_n43_8# 0.09fF
C465 enable_2/and_6/w_26_9# vdd 0.03fF
C466 vdd comparator_0/b2bar 1.10fF
C467 4bitadder_0/fulladder_3/XOR_1/w_n34_n1# vdd 0.02fF
C468 s0 decoder_0/and_1/w_n43_8# 0.09fF
C469 4bitadder_1/XOR_2/out 4bitadder_1/XOR_2/w_62_37# 0.02fF
C470 vdd decoder_0/and_2/w_26_9# 0.03fF
C471 4bitadder_0/fulladder_1/XOR_0/bbar 4bitadder_0/XOR_1/out 0.02fF
C472 4bitadder_0/XOR_3/bbar s0 0.02fF
C473 4bitadder_0/XOR_2/w_16_n1# vdd 0.02fF
C474 b0out_0 4bitadder_0/XOR_0/w_62_37# 0.02fF
C475 enable_0/and_4/w_26_9# vdd 0.03fF
C476 4bitadder_0/XOR_3/w_62_n20# 4bitadder_0/XOR_3/bbar 0.13fF
C477 enable_2/and_5/w_n43_8# enable_2/en 0.09fF
C478 vdd comparator_0/3input_AND_1/not_0/w_n2_10# 0.18fF
C479 4bitadder_1/fulladder_0/or_0/a_n15_32# 4bitadder_1/fulladder_0/or_0/w_n48_101# 0.05fF
C480 comparator_0/t3 comparator_0/t2 0.19fF
C481 enable_2/and_0/w_26_9# enable_2/and_0/a_n26_14# 0.09fF
C482 4bitadder_1/fulladder_0/XOR_1/bbar 4bitadder_1/fulladder_0/XOR_1/w_16_n1# 0.03fF
C483 AND_Block_0/and_0/w_n43_8# b0out_3 0.09fF
C484 comparator_0/4input_OR_1/y comparator_0/t2 0.18fF
C485 enable_1/en a0 0.24fF
C486 4bitadder_0/fulladder_0/axorb 4bitadder_0/fulladder_0/XOR_1/abar 0.13fF
C487 enable_1/and_6/w_26_9# b2out_1 0.03fF
C488 decoder_0/and_0/a_n26_14# decoder_0/and_0/w_26_9# 0.09fF
C489 4bitadder_1/fulladder_2/XOR_1/w_62_37# s2_sub 0.02fF
C490 s0 decoder_0/and_2/a 0.12fF
C491 comparator_0/xnor_3/not_0/in gnd 0.03fF
C492 4bitadder_0/fulladder_1/XOR_1/w_16_n1# 4bitadder_0/fulladder_1/XOR_1/bbar 0.03fF
C493 4bitadder_0/fulladder_1/XOR_1/w_62_n20# s1_add 0.04fF
C494 4bitadder_0/fulladder_1/XOR_1/w_n34_n1# 4bitadder_0/fulladder_1/XOR_1/abar 0.03fF
C495 enable_3/and_1/w_n43_8# vdd 0.07fF
C496 4bitadder_1/fulladder_1/XOR_0/w_n34_n1# 4bitadder_1/fulladder_1/XOR_0/abar 0.03fF
C497 comparator_0/and_1/w_26_9# comparator_0/and_1/a_n26_14# 0.09fF
C498 enable_3/and_6/a_n26_14# enable_3/and_6/w_26_9# 0.09fF
C499 enable_2/and_0/w_26_9# vdd 0.03fF
C500 comparator_0/xnor_1/XOR_0/w_62_37# a2out_2 0.02fF
C501 4bitadder_1/fulladder_1/and_0/a_n26_14# 4bitadder_1/c1 0.10fF
C502 4bitadder_0/fulladder_3/and_1/w_n43_8# a3out_0 0.09fF
C503 vdd 4bitadder_1/fulladder_1/XOR_0/w_n34_n1# 0.02fF
C504 boout_2 comparator_0/a3xnorb3 0.48fF
C505 enable_3/and_2/w_n43_8# a2 0.09fF
C506 vdd decoder_0/and_0/w_n43_8# 0.07fF
C507 4bitadder_1/c1 4bitadder_1/fulladder_1/XOR_1/w_16_n1# 0.11fF
C508 4bitadder_0/fulladder_0/XOR_1/w_n34_n1# vdd 0.02fF
C509 AND_Block_0/and_1/w_26_9# vdd 0.03fF
C510 b3out_0 s0 0.51fF
C511 AND_Block_0/and_2/w_n43_8# AND_Block_0/and_2/a_n26_14# 0.02fF
C512 vdd comparator_0/xnor_3/XOR_0/w_16_n1# 0.02fF
C513 comparator_0/xnor_1/XOR_0/w_62_n20# comparator_0/xnor_1/XOR_0/bbar 0.13fF
C514 enable_3/and_4/w_26_9# vdd 0.03fF
C515 4bitadder_1/c1 4bitadder_1/fulladder_1/XOR_1/abar 0.27fF
C516 4bitadder_1/fulladder_3/XOR_0/w_n34_n1# a3out_1 0.11fF
C517 4bitadder_1/fulladder_3/XOR_0/w_16_n1# 4bitadder_1/XOR_3/out 0.11fF
C518 enable_3/en enable_3/and_4/w_n43_8# 0.09fF
C519 vdd 4bitadder_1/c2 0.17fF
C520 4bitadder_1/b0xorM s0 0.26fF
C521 gnd 4bitadder_1/fulladder_3/or_0/a 0.01fF
C522 enable_3/and_5/w_n43_8# vdd 0.07fF
C523 4bitadder_1/fulladder_0/and_1/w_n43_8# 4bitadder_1/fulladder_0/and_1/a_n26_14# 0.02fF
C524 4bitadder_0/XOR_2/out 4bitadder_0/XOR_2/w_62_37# 0.02fF
C525 comparator_0/b1bar gnd 0.14fF
C526 enable_0/and_0/a_n26_14# a0 0.31fF
C527 4bitadder_1/fulladder_3/XOR_0/abar 4bitadder_1/XOR_3/out 0.25fF
C528 comparator_0/5input_AND_0/not_0/in comparator_0/5input_AND_0/w_n4_n20# 0.03fF
C529 4bitadder_0/fulladder_1/and_0/w_n43_8# vdd 0.07fF
C530 vdd comparator_0/not_5/w_n2_10# 0.18fF
C531 b1 vdd 0.47fF
C532 4bitadder_0/XOR_2/w_16_n1# s0 0.11fF
C533 4bitadder_0/fulladder_0/and_0/w_26_9# vdd 0.03fF
C534 comparator_0/a1xnorb1 boout_2 0.85fF
C535 4bitadder_0/fulladder_3/and_1/w_n43_8# vdd 0.07fF
C536 enable_0/and_7/w_26_9# b3out_0 0.03fF
C537 b1 a3 0.28fF
C538 comparator_0/not_2/w_n2_10# comparator_0/b2bar 0.03fF
C539 comparator_0/not_0/w_n2_10# comparator_0/b0bar 0.03fF
C540 4bitadder_0/fulladder_2/XOR_1/w_62_37# s2_add 0.02fF
C541 a2out_1 a3out_1 11.02fF
C542 enable_1/en enable_1/and_4/w_n43_8# 0.09fF
C543 4bitadder_1/XOR_3/out 4bitadder_1/XOR_3/w_62_37# 0.02fF
C544 comparator_0/3input_AND_1/w_n14_24# comparator_0/a2bar 0.16fF
C545 4bitadder_0/fulladder_2/or_0/a vdd 0.14fF
C546 4bitadder_0/fulladder_1/XOR_0/abar gnd 0.15fF
C547 4bitadder_0/fulladder_1/XOR_0/w_62_n20# 4bitadder_0/fulladder_1/XOR_0/abar 0.02fF
C548 4bitadder_0/XOR_2/abar s0 0.28fF
C549 enable_0/and_3/w_n43_8# vdd 0.07fF
C550 a0 gnd 0.27fF
C551 4bitadder_1/fulladder_3/XOR_1/w_62_n20# 4bitadder_1/fulladder_3/XOR_1/bbar 0.13fF
C552 4bitadder_0/XOR_0/abar s0 1.07fF
C553 4bitadder_0/c3 gnd 0.91fF
C554 a3out_2 b3out_2 3.20fF
C555 comparator_0/xnor_0/XOR_0/w_16_n1# comparator_0/xnor_0/XOR_0/bbar 0.03fF
C556 comparator_0/xnor_0/XOR_0/w_62_n20# comparator_0/xnor_0/not_0/in 0.04fF
C557 comparator_0/xnor_0/XOR_0/w_n34_n1# comparator_0/xnor_0/XOR_0/abar 0.03fF
C558 4bitadder_0/XOR_1/out s0 0.15fF
C559 s0 4bitadder_1/XOR_3/w_62_37# 0.13fF
C560 gnd 4bitadder_1/fulladder_1/or_0/a 0.01fF
C561 comparator_0/a2bar comparator_0/a3xnorb3 0.19fF
C562 enable_0/and_3/w_n43_8# a3 0.09fF
C563 4bitadder_1/c1 gnd 0.77fF
C564 vdd comparator_0/3input_AND_1/w_n14_24# 0.03fF
C565 decoder_0/and_2/w_26_9# decoder_0/and_2/a_n26_14# 0.09fF
C566 4bitadder_1/fulladder_2/or_0/a_n15_32# 4bitadder_1/fulladder_2/or_0/w_58_101# 0.13fF
C567 vdd comparator_0/5input_AND_0/w_106_n113# 0.04fF
C568 enable_3/en gnd 0.13fF
C569 vdd 4bitadder_1/XOR_2/w_n34_n1# 0.02fF
C570 b2out_1 4bitadder_1/XOR_2/abar 0.13fF
C571 a0 enable_3/and_0/a_n26_14# 0.31fF
C572 4bitadder_1/XOR_0/bbar 4bitadder_1/XOR_0/w_16_n1# 0.03fF
C573 vdd comparator_0/4input_AND_1/w_n8_2# 0.02fF
C574 vdd s3_sub 0.10fF
C575 4bitadder_1/XOR_1/out 4bitadder_1/fulladder_1/XOR_0/abar 0.25fF
C576 enable_2/and_6/a_n26_14# b2 0.31fF
C577 comparator_0/t8 comparator_0/t5 0.21fF
C578 vdd comparator_0/a3xnorb3 1.70fF
C579 4bitadder_0/fulladder_3/XOR_0/w_n34_n1# a3out_0 0.11fF
C580 4bitadder_0/fulladder_3/XOR_0/w_16_n1# 4bitadder_0/XOR_3/out 0.11fF
C581 AND_Block_0/and_3/w_n43_8# AND_Block_0/and_3/a_n26_14# 0.02fF
C582 comparator_0/4input_AND_0/not_0/in comparator_0/4input_AND_0/w_n47_52# 0.02fF
C583 comparator_0/b1bar comparator_0/a2xnorb2 0.51fF
C584 4bitadder_0/fulladder_3/axorb vdd 0.15fF
C585 4bitadder_0/fulladder_0/XOR_1/bbar s0 0.02fF
C586 4bitadder_0/fulladder_0/and_1/w_n43_8# a0out_0 0.09fF
C587 4bitadder_0/fulladder_0/and_1/w_n43_8# vdd 0.07fF
C588 enable_3/and_7/w_n43_8# enable_3/en 0.09fF
C589 enable_2/and_7/w_n43_8# enable_2/en 0.09fF
C590 b1out_2 gnd 1.06fF
C591 a3out_2 a1out_2 0.75fF
C592 enable_1/en a2 0.28fF
C593 a0_out1 gnd 0.56fF
C594 4bitadder_1/fulladder_0/XOR_1/w_62_37# 4bitadder_1/fulladder_0/axorb 0.02fF
C595 comparator_0/a3bar comparator_0/and_1/w_n43_8# 0.09fF
C596 4bitadder_1/b0xorM 4bitadder_1/XOR_0/w_62_n20# 0.04fF
C597 vdd 4bitadder_1/fulladder_0/and_0/w_n43_8# 0.07fF
C598 4bitadder_0/fulladder_3/XOR_0/abar 4bitadder_0/XOR_3/out 0.25fF
C599 AND_Block_0/and_1/w_26_9# out1 0.03fF
C600 enable_3/and_3/w_n43_8# vdd 0.07fF
C601 4bitadder_1/fulladder_0/and_0/w_n43_8# 4bitadder_1/fulladder_0/axorb 0.09fF
C602 vdd comparator_0/4input_AND_2/not_0/w_n2_10# 0.18fF
C603 4bitadder_1/c1 4bitadder_1/fulladder_0/or_0/w_58_101# 0.02fF
C604 4bitadder_0/fulladder_1/or_0/w_n48_101# vdd 0.05fF
C605 vdd 4bitadder_1/fulladder_0/or_0/a 0.14fF
C606 vdd comparator_0/xnor_2/XOR_0/w_n34_n1# 0.02fF
C607 enable_3/and_3/w_n43_8# a3 0.09fF
C608 a1out_3 vdd 0.16fF
C609 4bitadder_1/c2 4bitadder_1/fulladder_2/XOR_1/bbar 0.02fF
C610 b2out_2 boout_2 0.30fF
C611 boout_2 comparator_0/5input_AND_1/w_n4_n20# 0.18fF
C612 4bitadder_0/fulladder_1/and_0/a_n26_14# 4bitadder_0/c1 0.10fF
C613 a2out_0 a3out_0 1.82fF
C614 enable_3/en decoder_0/and_3/w_26_9# 0.03fF
C615 vdd comparator_0/4input_AND_2/w_29_n46# 0.02fF
C616 enable_2/and_5/a_n26_14# b1 0.31fF
C617 4bitadder_0/XOR_3/out 4bitadder_0/XOR_3/w_62_37# 0.02fF
C618 4bitadder_0/fulladder_3/XOR_1/w_62_n20# 4bitadder_0/fulladder_3/XOR_1/bbar 0.13fF
C619 4bitadder_0/fulladder_1/axorb 4bitadder_0/fulladder_1/XOR_1/abar 0.13fF
C620 4bitadder_0/fulladder_0/or_0/a_n15_32# 4bitadder_0/fulladder_0/or_0/b 0.19fF
C621 enable_0/and_1/w_26_9# a1out_0 0.03fF
C622 vdd 4bitadder_1/fulladder_0/XOR_0/w_16_n1# 0.02fF
C623 4bitadder_1/fulladder_0/and_0/w_26_9# 4bitadder_1/fulladder_0/and_0/a_n26_14# 0.09fF
C624 vdd comparator_0/a1xnorb1 0.87fF
C625 comparator_0/4input_AND_1/not_0/in comparator_0/4input_AND_1/not_0/w_n2_10# 0.09fF
C626 comparator_0/xnor_2/XOR_0/w_62_37# b1out_2 0.13fF
C627 vdd comparator_0/not_1/w_n2_10# 0.18fF
C628 4bitadder_0/fulladder_3/XOR_0/w_n34_n1# vdd 0.02fF
C629 gnd a3out_1 1.05fF
C630 4bitadder_1/fulladder_1/and_1/w_n43_8# a1out_1 0.09fF
C631 b1out_2 comparator_0/4input_AND_2/w_n8_2# 0.16fF
C632 enable_2/and_0/w_n43_8# enable_2/and_0/a_n26_14# 0.02fF
C633 enable_0/and_1/a_n26_14# a1 0.31fF
C634 b1out_2 comparator_0/xnor_2/not_0/in 0.13fF
C635 a1out_2 comparator_0/xnor_2/XOR_0/abar 0.13fF
C636 4bitadder_0/XOR_0/bbar 4bitadder_0/XOR_0/w_16_n1# 0.03fF
C637 4bitadder_0/fulladder_2/or_0/a_n15_32# 4bitadder_0/fulladder_2/or_0/b 0.19fF
C638 enable_1/en enable_1/and_7/w_n43_8# 0.09fF
C639 a0_out1 4bitadder_1/fulladder_0/XOR_0/w_62_37# 0.02fF
C640 AND_Block_0/and_2/w_26_9# out2 0.03fF
C641 b1out_2 comparator_0/a2xnorb2 0.26fF
C642 enable_2/en gnd 0.16fF
C643 enable_0/and_6/w_26_9# b2out_0 0.03fF
C644 4bitadder_1/fulladder_2/and_1/w_n43_8# 4bitadder_1/fulladder_2/and_1/a_n26_14# 0.02fF
C645 enable_2/and_0/w_n43_8# vdd 0.07fF
C646 enable_1/and_6/w_n43_8# b2 0.09fF
C647 4bitadder_1/XOR_1/out s0 0.15fF
C648 4bitadder_1/fulladder_0/XOR_1/w_62_37# s0 0.13fF
C649 s0 4bitadder_1/XOR_2/bbar 0.02fF
C650 a2out_0 vdd 0.35fF
C651 enable_2/and_1/w_26_9# enable_2/and_1/a_n26_14# 0.09fF
C652 gnd 4bitadder_1/fulladder_2/XOR_1/abar 0.15fF
C653 a2out_2 gnd 0.88fF
C654 a2 gnd 0.27fF
C655 4bitadder_1/fulladder_1/axorb 4bitadder_1/fulladder_1/XOR_0/w_62_37# 0.02fF
C656 enable_2/and_1/w_n43_8# a1 0.09fF
C657 decoder_0/and_1/a_n26_14# decoder_0/and_1/w_n43_8# 0.02fF
C658 4bitadder_1/fulladder_3/and_0/a_n26_14# 4bitadder_1/fulladder_3/and_0/w_26_9# 0.09fF
C659 4bitadder_1/fulladder_0/and_0/w_n43_8# s0 0.09fF
C660 4bitadder_0/fulladder_0/XOR_0/w_n34_n1# vdd 0.02fF
C661 4bitadder_0/fulladder_0/XOR_0/w_n34_n1# a0out_0 0.11fF
C662 4bitadder_0/fulladder_0/XOR_0/w_16_n1# 4bitadder_0/b0xorM 0.11fF
C663 enable_0/and_4/w_n43_8# b0 0.09fF
C664 b2out_2 comparator_0/a2bar 0.27fF
C665 a1out_1 b2out_1 0.25fF
C666 4bitadder_0/c2 4bitadder_0/fulladder_2/XOR_1/bbar 0.02fF
C667 enable_3/and_7/a_n26_14# enable_3/and_7/w_n43_8# 0.02fF
C668 comparator_0/5input_AND_1/not_0/in comparator_0/5input_AND_1/w_106_n113# 0.03fF
C669 4bitadder_0/fulladder_1/XOR_1/w_16_n1# vdd 0.02fF
C670 enable_2/and_2/w_26_9# vdd 0.03fF
C671 comparator_0/a0xnorb0 comparator_0/xnor_3/not_0/w_n2_10# 0.03fF
C672 vdd 4bitadder_1/fulladder_3/and_0/w_26_9# 0.03fF
C673 a1 enable_3/and_1/a_n26_14# 0.31fF
C674 4bitadder_1/XOR_0/w_62_37# b0out_1 0.02fF
C675 4bitadder_0/fulladder_0/XOR_0/abar 4bitadder_0/b0xorM 0.25fF
C676 4bitadder_1/fulladder_1/and_0/w_26_9# 4bitadder_1/fulladder_1/or_0/a 0.03fF
C677 4bitadder_0/c1 4bitadder_0/XOR_1/out 0.37fF
C678 enable_2/and_0/w_26_9# a0out_2 0.03fF
C679 a1out_1 4bitadder_1/fulladder_1/and_1/a_n26_14# 0.10fF
C680 enable_1/and_5/a_n26_14# enable_1/and_5/w_26_9# 0.09fF
C681 vdd b2out_2 1.44fF
C682 vdd comparator_0/5input_AND_1/w_n4_n20# 0.05fF
C683 enable_1/en b0 0.28fF
C684 enable_0/en a0 0.38fF
C685 comparator_0/4input_AND_0/not_0/in gnd 0.03fF
C686 comparator_0/a0bar comparator_0/not_4/w_n2_10# 0.03fF
C687 4bitadder_0/fulladder_2/or_0/w_58_101# vdd 0.05fF
C688 enable_2/and_4/w_26_9# boout_2 0.03fF
C689 enable_1/and_5/w_n43_8# b1 0.09fF
C690 b2out_3 b1out_3 29.73fF
C691 4bitadder_1/fulladder_0/and_1/w_26_9# 4bitadder_1/fulladder_0/or_0/b 0.03fF
C692 comparator_0/4input_OR_0/y comparator_0/t5 0.18fF
C693 4bitadder_0/fulladder_0/XOR_1/w_62_n20# 4bitadder_0/fulladder_0/XOR_1/bbar 0.13fF
C694 b0out_0 a3out_0 0.12fF
C695 comparator_0/4input_AND_1/not_0/in gnd 0.21fF
C696 decoder_0/and_2/a s1 0.24fF
C697 4bitadder_1/fulladder_1/axorb 4bitadder_1/fulladder_1/XOR_1/abar 0.13fF
C698 boout_2 comparator_0/xnor_3/not_0/in 0.13fF
C699 a0out_2 comparator_0/xnor_3/XOR_0/abar 0.13fF
C700 comparator_0/not_0/w_n2_10# boout_2 0.09fF
C701 4bitadder_0/fulladder_2/and_1/w_n43_8# 4bitadder_0/fulladder_2/and_1/a_n26_14# 0.02fF
C702 enable_3/and_4/w_n43_8# b0 0.09fF
C703 b3out_2 enable_2/and_7/w_26_9# 0.03fF
C704 a2out_2 comparator_0/a2xnorb2 0.17fF
C705 comparator_0/4input_AND_1/not_0/in comparator_0/4input_AND_1/w_n47_52# 0.02fF
C706 a3out_1 4bitadder_1/fulladder_3/and_1/a_n26_14# 0.10fF
C707 enable_3/and_6/w_26_9# b2out_3 0.03fF
C708 a2out_0 s0 0.31fF
C709 4bitadder_1/c2 4bitadder_1/fulladder_2/axorb 0.54fF
C710 4bitadder_0/fulladder_3/and_0/a_n26_14# 4bitadder_0/fulladder_3/and_0/w_26_9# 0.09fF
C711 vdd s0_sub 0.19fF
C712 4bitadder_1/b0xorM 4bitadder_1/fulladder_0/XOR_0/bbar 0.02fF
C713 vdd enable_1/and_1/w_26_9# 0.03fF
C714 4bitadder_0/c1 4bitadder_0/fulladder_1/and_0/w_n43_8# 0.09fF
C715 4bitadder_1/fulladder_1/or_0/w_n48_101# 4bitadder_1/fulladder_1/or_0/a 0.12fF
C716 vdd comparator_0/3input_AND_0/w_69_n71# 0.03fF
C717 enable_1/and_3/w_26_9# vdd 0.03fF
C718 comparator_0/and_0/w_n43_8# comparator_0/and_0/a_n26_14# 0.02fF
C719 comparator_0/and_0/w_26_9# comparator_0/t5 0.03fF
C720 s0 4bitadder_1/XOR_1/abar 0.25fF
C721 4bitadder_0/fulladder_1/or_0/b gnd 0.37fF
C722 enable_3/and_4/w_26_9# b0out_3 0.03fF
C723 vdd comparator_0/t7 0.04fF
C724 4bitadder_0/fulladder_0/axorb 4bitadder_0/fulladder_0/XOR_1/w_62_37# 0.02fF
C725 enable_0/and_2/a_n26_14# a2 0.31fF
C726 b2out_3 gnd 0.24fF
C727 4bitadder_1/fulladder_2/XOR_0/abar a2out_1 0.13fF
C728 a2out_1 b2out_1 0.16fF
C729 b3out_2 comparator_0/and_1/a_n26_14# 0.10fF
C730 4bitadder_1/c3 a3out_1 0.40fF
C731 comparator_0/4input_AND_0/not_0/in comparator_0/a2xnorb2 0.18fF
C732 b0out_0 vdd 0.13fF
C733 enable_2/en enable_2/and_2/w_n43_8# 0.09fF
C734 4bitadder_0/fulladder_1/and_1/w_26_9# vdd 0.03fF
C735 enable_2/and_1/w_n43_8# vdd 0.07fF
C736 a0 a1 0.31fF
C737 4bitadder_1/XOR_0/w_62_37# s0 0.13fF
C738 4bitadder_1/fulladder_1/axorb gnd 0.09fF
C739 enable_2/and_2/w_26_9# enable_2/and_2/a_n26_14# 0.09fF
C740 b2out_3 a3out_3 0.13fF
C741 b0 gnd 0.30fF
C742 comparator_0/t7 comparator_0/t6 0.27fF
C743 comparator_0/4input_AND_1/not_0/in comparator_0/a2xnorb2 0.18fF
C744 enable_2/and_2/w_n43_8# a2 0.09fF
C745 4bitadder_1/fulladder_2/XOR_1/w_62_n20# 4bitadder_1/fulladder_2/XOR_1/abar 0.02fF
C746 4bitadder_0/XOR_0/w_16_n1# vdd 0.02fF
C747 enable_3/and_7/w_26_9# vdd 0.03fF
C748 enable_1/and_1/a_n26_14# enable_1/and_1/w_26_9# 0.09fF
C749 a0out_2 comparator_0/a3xnorb3 0.28fF
C750 comparator_0/not_2/w_n2_10# b2out_2 0.09fF
C751 enable_2/and_1/w_26_9# a1out_2 0.03fF
C752 4bitadder_1/c1 4bitadder_1/fulladder_1/XOR_1/w_62_37# 0.13fF
C753 AND_Block_0/and_0/a_n26_14# AND_Block_0/and_0/w_26_9# 0.09fF
C754 vdd 4bitadder_1/fulladder_1/XOR_1/w_n34_n1# 0.02fF
C755 b3out_0 4bitadder_0/XOR_3/w_n34_n1# 0.11fF
C756 enable_1/and_2/w_26_9# enable_1/and_2/a_n26_14# 0.09fF
C757 b3 a0 0.32fF
C758 enable_3/en a1 0.25fF
C759 a0out_3 gnd 0.11fF
C760 enable_2/and_4/w_26_9# vdd 0.03fF
C761 a3out_0 4bitadder_0/fulladder_3/and_1/a_n26_14# 0.10fF
C762 a2 enable_3/and_2/a_n26_14# 0.31fF
C763 4bitadder_1/c1 s1_sub 0.04fF
C764 4bitadder_0/c2 4bitadder_0/fulladder_2/axorb 0.54fF
C765 4bitadder_1/fulladder_3/XOR_0/w_62_37# 4bitadder_1/XOR_3/out 0.13fF
C766 comparator_0/not_0/w_n2_10# vdd 0.18fF
C767 b1out_1 4bitadder_1/XOR_1/abar 0.13fF
C768 4bitadder_0/XOR_3/out gnd 0.42fF
C769 a2out_0 b1out_0 0.14fF
C770 s0_sub s0 0.04fF
C771 enable_3/en b3 0.32fF
C772 enable_1/and_0/w_n43_8# a0 0.09fF
C773 enable_0/en a2 0.38fF
C774 vdd 4bitadder_1/fulladder_2/and_0/w_n43_8# 0.07fF
C775 4bitadder_0/fulladder_0/axorb gnd 0.09fF
C776 enable_2/and_7/a_n26_14# enable_2/and_7/w_26_9# 0.09fF
C777 b1out_2 boout_2 0.73fF
C778 4bitadder_0/XOR_1/out 4bitadder_0/XOR_1/w_62_n20# 0.04fF
C779 4bitadder_0/fulladder_2/XOR_0/abar a2out_0 0.13fF
C780 enable_0/en decoder_0/and_0/w_26_9# 0.03fF
C781 4bitadder_1/XOR_1/w_62_37# s0 0.13fF
C782 comparator_0/a1xnorb1 a0out_2 0.40fF
C783 4bitadder_0/XOR_2/w_62_37# s0 0.13fF
C784 4bitadder_0/c3 a3out_0 0.36fF
C785 enable_0/and_7/w_n43_8# enable_0/and_7/a_n26_14# 0.02fF
C786 enable_1/and_2/w_n43_8# vdd 0.07fF
C787 comparator_0/xnor_3/XOR_0/w_62_37# comparator_0/xnor_3/not_0/in 0.02fF
C788 4bitadder_0/fulladder_1/XOR_0/w_16_n1# 4bitadder_0/fulladder_1/XOR_0/bbar 0.03fF
C789 4bitadder_0/fulladder_1/XOR_0/w_n34_n1# 4bitadder_0/fulladder_1/XOR_0/abar 0.03fF
C790 b0out_0 s0 0.15fF
C791 a2out_2 comparator_0/3input_AND_0/w_32_n21# 0.16fF
C792 b3out_2 gnd 0.98fF
C793 vdd 4bitadder_1/fulladder_3/or_0/a 0.14fF
C794 gnd 4bitadder_1/fulladder_2/XOR_0/abar 0.15fF
C795 comparator_0/xnor_0/XOR_0/w_16_n1# b3out_2 0.11fF
C796 gnd b2out_1 0.92fF
C797 vdd comparator_0/5input_AND_0/not_0/w_n2_10# 0.17fF
C798 4bitadder_1/XOR_2/out s0 0.19fF
C799 comparator_0/b1bar vdd 0.20fF
C800 4bitadder_0/fulladder_2/XOR_1/w_62_n20# 4bitadder_0/fulladder_2/XOR_1/abar 0.02fF
C801 4bitadder_1/XOR_2/w_62_37# b2out_1 0.02fF
C802 4bitadder_1/fulladder_3/axorb 4bitadder_1/fulladder_3/XOR_0/w_62_n20# 0.04fF
C803 a1out_3 b0out_3 0.21fF
C804 comparator_0/3input_AND_1/w_69_n71# comparator_0/a3xnorb3 0.16fF
C805 enable_0/en enable_0/and_5/w_n43_8# 0.09fF
C806 a3out_1 b3out_1 0.20fF
C807 a0_out1 4bitadder_1/fulladder_0/XOR_0/w_n34_n1# 0.11fF
C808 comparator_0/4input_OR_0/w_n58_n43# comparator_0/t7 0.13fF
C809 enable_2/and_0/a_n26_14# a0 0.31fF
C810 b3out_2 comparator_0/xnor_0/XOR_0/abar 0.30fF
C811 4bitadder_0/XOR_0/w_16_n1# s0 0.11fF
C812 4bitadder_0/fulladder_1/XOR_0/w_16_n1# vdd 0.02fF
C813 4bitadder_0/b0xorM gnd 0.42fF
C814 vdd comparator_0/5input_AND_0/w_31_n55# 0.06fF
C815 vdd comparator_0/xnor_0/XOR_0/w_n34_n1# 0.02fF
C816 4bitadder_1/XOR_2/w_62_n20# 4bitadder_1/XOR_2/bbar 0.13fF
C817 4bitadder_1/fulladder_2/and_0/w_26_9# 4bitadder_1/fulladder_2/or_0/a 0.03fF
C818 enable_0/and_3/a_n26_14# a3 0.31fF
C819 a3out_0 a0_out1 0.21fF
C820 comparator_0/a1bar comparator_0/not_5/w_n2_10# 0.03fF
C821 comparator_0/t4 comparator_0/5input_AND_1/not_0/w_n2_10# 0.03fF
C822 b3out_2 comparator_0/not_3/w_n2_10# 0.09fF
C823 comparator_0/xnor_0/not_0/w_n2_10# comparator_0/a3xnorb3 0.03fF
C824 4bitadder_0/fulladder_3/XOR_0/w_62_37# 4bitadder_0/XOR_3/out 0.13fF
C825 enable_2/en a1 0.28fF
C826 AND_Block_0/and_3/w_n43_8# a3out_3 0.09fF
C827 a0 vdd 0.41fF
C828 b3out_2 comparator_0/and_1/w_n43_8# 0.09fF
C829 4bitadder_0/c3 vdd 0.12fF
C830 4bitadder_0/b0xorM 4bitadder_0/XOR_0/w_62_37# 0.02fF
C831 a1out_2 gnd 0.83fF
C832 enable_2/and_7/w_n43_8# enable_2/and_7/a_n26_14# 0.02fF
C833 vdd comparator_0/a3bar 0.04fF
C834 enable_2/en enable_2/and_4/w_n43_8# 0.09fF
C835 vdd 4bitadder_1/XOR_1/w_n34_n1# 0.02fF
C836 comparator_0/t5 gnd 0.34fF
C837 comparator_0/4input_OR_1/y gnd 0.03fF
C838 a3out_2 comparator_0/b3bar 3.31fF
C839 enable_2/and_3/w_n43_8# vdd 0.07fF
C840 vdd 4bitadder_1/fulladder_1/or_0/a 0.14fF
C841 a1out_2 comparator_0/4input_AND_1/w_n47_52# 0.16fF
C842 vdd 4bitadder_1/c1 0.12fF
C843 4bitadder_1/XOR_1/w_62_37# b1out_1 0.02fF
C844 comparator_0/4input_AND_2/not_0/in comparator_0/a3xnorb3 0.18fF
C845 a0 a3 0.31fF
C846 a1 a2 0.40fF
C847 enable_2/and_3/w_26_9# enable_2/and_3/a_n26_14# 0.09fF
C848 a0out_0 4bitadder_0/fulladder_0/and_1/a_n26_14# 0.10fF
C849 vdd comparator_0/and_1/w_26_9# 0.03fF
C850 enable_2/en b3 0.22fF
C851 enable_2/and_3/w_n43_8# a3 0.09fF
C852 comparator_0/4input_OR_1/w_n58_n43# comparator_0/t4 0.13fF
C853 4bitadder_0/fulladder_1/axorb 4bitadder_0/fulladder_1/XOR_1/w_62_37# 0.02fF
C854 4bitadder_0/c1 4bitadder_0/fulladder_1/XOR_1/w_16_n1# 0.11fF
C855 4bitadder_0/fulladder_0/or_0/w_58_101# vdd 0.05fF
C856 enable_3/en vdd 0.68fF
C857 vdd decoder_0/and_3/w_n43_8# 0.07fF
C858 decoder_0/and_0/w_n43_8# decoder_0/and_2/a 0.09fF
C859 comparator_0/3input_AND_0/not_0/in comparator_0/a3xnorb3 0.19fF
C860 a2out_2 boout_2 0.51fF
C861 b2out_2 a0out_2 0.42fF
C862 vdd comparator_0/4input_AND_2/w_n47_52# 0.02fF
C863 enable_1/and_3/w_26_9# enable_1/and_3/a_n26_14# 0.09fF
C864 b3 a2 0.31fF
C865 4bitadder_1/fulladder_3/XOR_0/w_62_n20# 4bitadder_1/fulladder_3/XOR_0/bbar 0.13fF
C866 comparator_0/a0xnorb0 gnd 0.36fF
C867 comparator_0/4input_AND_2/not_0/w_n2_10# comparator_0/4input_AND_2/not_0/in 0.09fF
C868 enable_3/en a3 0.23fF
C869 enable_3/and_7/a_n26_14# b3 0.31fF
C870 4bitadder_0/fulladder_0/or_0/w_n48_101# 4bitadder_0/fulladder_0/or_0/b 0.12fF
C871 vdd b1out_2 1.29fF
C872 4bitadder_0/c1 4bitadder_0/fulladder_1/XOR_1/abar 0.27fF
C873 4bitadder_1/fulladder_2/and_0/a_n26_14# 4bitadder_1/c2 0.10fF
C874 vdd a0_out1 0.26fF
C875 a3 enable_3/and_3/a_n26_14# 0.31fF
C876 comparator_0/xnor_2/XOR_0/w_62_37# a1out_2 0.02fF
C877 4bitadder_1/fulladder_0/XOR_0/bbar 4bitadder_1/fulladder_0/XOR_0/w_16_n1# 0.03fF
C878 vdd 4bitadder_1/fulladder_0/or_0/w_n48_101# 0.05fF
C879 4bitadder_0/fulladder_3/axorb 4bitadder_0/fulladder_3/XOR_0/w_62_n20# 0.04fF
C880 4bitadder_0/fulladder_1/and_0/a_n26_14# 4bitadder_0/fulladder_1/and_0/w_n43_8# 0.02fF
C881 comparator_0/a1bar comparator_0/a3xnorb3 0.36fF
C882 comparator_0/4input_AND_2/not_0/in comparator_0/4input_AND_2/w_29_n46# 0.02fF
C883 decoder_0/and_3/w_26_9# decoder_0/and_3/a_n26_14# 0.09fF
C884 4bitadder_0/fulladder_1/or_0/w_58_101# 4bitadder_0/c2 0.02fF
C885 comparator_0/4input_OR_1/w_n58_n43# comparator_0/t3 0.13fF
C886 4bitadder_0/fulladder_1/or_0/a gnd 0.01fF
C887 comparator_0/xnor_2/XOR_0/w_62_n20# comparator_0/xnor_2/XOR_0/bbar 0.13fF
C888 4bitadder_0/XOR_1/bbar s0 0.02fF
C889 4bitadder_0/fulladder_0/axorb 4bitadder_0/fulladder_0/XOR_0/w_62_37# 0.02fF
C890 enable_0/en b0 0.38fF
C891 4bitadder_0/XOR_2/w_62_n20# 4bitadder_0/XOR_2/bbar 0.13fF
C892 enable_1/and_7/a_n26_14# enable_1/and_7/w_n43_8# 0.02fF
C893 vdd comparator_0/3input_AND_0/not_0/w_n2_10# 0.18fF
C894 4bitadder_0/fulladder_2/and_0/w_26_9# 4bitadder_0/fulladder_2/or_0/a 0.03fF
C895 comparator_0/4input_OR_1/y comparator_0/4input_OR_1/w_n58_n43# 0.02fF
C896 4bitadder_1/XOR_0/bbar s0 0.02fF
C897 a1out_2 comparator_0/a2xnorb2 0.61fF
C898 enable_0/and_6/w_n43_8# enable_0/and_6/a_n26_14# 0.02fF
C899 a3out_1 b0out_1 0.13fF
C900 4bitadder_1/fulladder_2/and_1/w_n43_8# 4bitadder_1/XOR_2/out 0.09fF
C901 enable_1/and_1/w_n43_8# enable_1/en 0.09fF
C902 AND_Block_0/and_1/a_n26_14# AND_Block_0/and_1/w_26_9# 0.09fF
C903 4bitadder_0/XOR_3/abar gnd 0.20fF
C904 enable_1/and_4/w_n43_8# vdd 0.07fF
C905 4bitadder_0/fulladder_1/and_1/w_26_9# 4bitadder_0/fulladder_1/and_1/a_n26_14# 0.09fF
C906 out2 gnd 0.01fF
C907 4bitadder_1/XOR_1/w_16_n1# 4bitadder_1/XOR_1/bbar 0.03fF
C908 vdd a3out_1 0.15fF
C909 enable_1/and_6/w_n43_8# enable_1/en 0.09fF
C910 enable_1/and_5/w_n43_8# enable_1/and_5/a_n26_14# 0.02fF
C911 b3 enable_1/and_7/w_n43_8# 0.09fF
C912 comparator_0/t6 comparator_0/3input_AND_0/not_0/w_n2_10# 0.03fF
C913 enable_1/en b2 0.28fF
C914 4bitadder_1/fulladder_3/axorb 4bitadder_1/fulladder_3/XOR_1/w_n34_n1# 0.11fF
C915 4bitadder_0/fulladder_2/axorb gnd 0.09fF
C916 4bitadder_0/fulladder_0/XOR_0/w_62_37# 4bitadder_0/b0xorM 0.13fF
C917 comparator_0/a0xnorb0 comparator_0/a2xnorb2 0.36fF
C918 comparator_0/xnor_1/XOR_0/abar gnd 0.14fF
C919 comparator_0/5input_AND_1/not_0/in comparator_0/5input_AND_1/w_31_n55# 0.03fF
C920 enable_2/and_1/a_n26_14# a1 0.31fF
C921 4bitadder_0/fulladder_3/XOR_0/w_62_n20# 4bitadder_0/fulladder_3/XOR_0/bbar 0.13fF
C922 s0 decoder_0/and_3/w_n43_8# 0.09fF
C923 vdd 4bitadder_1/fulladder_2/XOR_1/w_16_n1# 0.02fF
C924 enable_2/en vdd 1.03fF
C925 4bitadder_0/fulladder_2/or_0/a_n15_32# 4bitadder_0/fulladder_2/or_0/w_58_101# 0.13fF
C926 enable_0/and_4/a_n26_14# b0 0.31fF
C927 s1_add vdd 0.19fF
C928 a0_out1 s0 0.29fF
C929 vdd a2out_2 1.48fF
C930 enable_2/en a3 0.28fF
C931 a2 vdd 0.41fF
C932 4bitadder_1/fulladder_2/axorb 4bitadder_1/XOR_2/out 0.13fF
C933 4bitadder_1/fulladder_1/axorb 4bitadder_1/fulladder_1/XOR_1/w_62_37# 0.02fF
C934 4bitadder_1/XOR_1/out 4bitadder_1/fulladder_1/XOR_0/w_16_n1# 0.11fF
C935 a1 b0 0.37fF
C936 a2 a3 0.31fF
C937 vdd 4bitadder_1/fulladder_3/or_0/w_58_101# 0.05fF
C938 enable_2/and_4/w_26_9# enable_2/and_4/a_n26_14# 0.09fF
C939 vdd decoder_0/and_0/w_26_9# 0.03fF
C940 enable_0/and_2/w_26_9# a2out_0 0.03fF
C941 enable_2/and_4/w_n43_8# b0 0.09fF
C942 comparator_0/xnor_3/XOR_0/w_62_n20# comparator_0/xnor_3/XOR_0/bbar 0.13fF
C943 4bitadder_1/XOR_1/w_n34_n1# b1out_1 0.11fF
C944 4bitadder_1/XOR_0/bbar 4bitadder_1/XOR_0/w_62_n20# 0.13fF
C945 comparator_0/3input_AND_1/not_0/in comparator_0/3input_AND_1/w_32_n21# 0.02fF
C946 4bitadder_0/fulladder_2/and_1/w_n43_8# 4bitadder_0/XOR_2/out 0.09fF
C947 4bitadder_1/XOR_3/out a3out_1 2.13fF
C948 4bitadder_1/fulladder_3/and_1/w_26_9# 4bitadder_1/fulladder_3/or_0/b 0.03fF
C949 enable_1/and_4/w_26_9# enable_1/and_4/a_n26_14# 0.09fF
C950 b3 b0 0.35fF
C951 vdd comparator_0/not_7/w_n2_10# 0.26fF
C952 comparator_0/4input_OR_1/NOT_0/w_n2_10# comparator_0/4input_OR_1/y 0.09fF
C953 4bitadder_0/XOR_1/w_16_n1# 4bitadder_0/XOR_1/bbar 0.03fF
C954 4bitadder_1/c1 4bitadder_1/fulladder_1/and_0/w_n43_8# 0.09fF
C955 4bitadder_0/fulladder_3/XOR_1/abar gnd 0.15fF
C956 comparator_0/b2bar comparator_0/a3xnorb3 0.38fF
C957 b0 enable_3/and_4/a_n26_14# 0.31fF
C958 b2out_3 AND_Block_0/and_2/w_n43_8# 0.09fF
C959 vdd enable_0/and_5/w_n43_8# 0.07fF
C960 4bitadder_0/fulladder_3/axorb 4bitadder_0/fulladder_3/XOR_1/w_n34_n1# 0.11fF
C961 enable_1/and_0/w_26_9# vdd 0.03fF
C962 4bitadder_1/fulladder_2/XOR_0/w_62_37# a2out_1 0.02fF
C963 vdd comparator_0/3input_AND_0/w_n14_24# 0.03fF
C964 4bitadder_1/fulladder_0/XOR_0/abar gnd 0.15fF
C965 b2 gnd 0.30fF
C966 4bitadder_1/fulladder_2/axorb 4bitadder_1/fulladder_2/and_0/w_n43_8# 0.09fF
C967 a1out_0 gnd 0.92fF
C968 enable_3/and_5/w_n43_8# b1 0.09fF
C969 vdd enable_1/and_7/w_n43_8# 0.07fF
C970 gnd 4bitadder_1/fulladder_2/or_0/b 0.37fF
C971 4bitadder_1/fulladder_2/XOR_0/bbar 4bitadder_1/XOR_2/out 0.02fF
C972 4bitadder_1/XOR_2/out 4bitadder_1/XOR_2/w_62_n20# 0.04fF
C973 AND_Block_0/and_0/w_n43_8# AND_Block_0/and_0/a_n26_14# 0.02fF
C974 4bitadder_1/b0xorM 4bitadder_1/fulladder_0/XOR_0/w_16_n1# 0.11fF
C975 enable_1/and_0/a_n26_14# enable_1/and_0/w_n43_8# 0.02fF
C976 enable_0/and_0/w_n43_8# enable_0/and_0/a_n26_14# 0.02fF
C977 4bitadder_0/fulladder_2/axorb 4bitadder_0/XOR_2/out 0.13fF
C978 comparator_0/3input_AND_0/not_0/in comparator_0/3input_AND_0/w_69_n71# 0.02fF
C979 vdd 4bitadder_1/fulladder_2/and_1/w_26_9# 0.03fF
C980 a2out_3 b2out_3 2.92fF
C981 4bitadder_0/fulladder_0/XOR_0/w_62_n20# 4bitadder_0/fulladder_0/XOR_0/bbar 0.13fF
C982 AND_Block_0/and_0/a_n26_14# b0out_3 0.31fF
C983 comparator_0/4input_OR_1/w_n58_n43# comparator_0/t2 0.13fF
C984 enable_3/and_6/w_n43_8# enable_3/and_6/a_n26_14# 0.02fF
C985 enable_2/and_6/w_n43_8# vdd 0.07fF
C986 4bitadder_1/fulladder_2/XOR_1/w_16_n1# 4bitadder_1/fulladder_2/XOR_1/bbar 0.03fF
C987 4bitadder_1/fulladder_2/XOR_1/w_62_n20# s2_sub 0.04fF
C988 4bitadder_1/fulladder_2/XOR_1/w_n34_n1# 4bitadder_1/fulladder_2/XOR_1/abar 0.03fF
C989 comparator_0/4input_OR_0/NOT_0/w_n2_10# comparator_0/4input_OR_0/y 0.09fF
C990 4bitadder_0/fulladder_1/axorb 4bitadder_0/fulladder_1/XOR_0/w_62_37# 0.02fF
C991 4bitadder_0/fulladder_0/XOR_1/abar gnd 0.15fF
C992 b2out_3 vdd 0.14fF
C993 b3out_2 boout_2 0.36fF
C994 b2out_0 4bitadder_0/XOR_2/w_n34_n1# 0.11fF
C995 4bitadder_0/XOR_0/bbar 4bitadder_0/XOR_0/w_62_n20# 0.13fF
C996 enable_2/and_2/a_n26_14# a2 0.31fF
C997 comparator_0/xnor_1/XOR_0/w_62_37# comparator_0/xnor_1/not_0/in 0.02fF
C998 4bitadder_0/fulladder_0/or_0/w_n48_101# 4bitadder_0/fulladder_0/or_0/a 0.12fF
C999 a3out_1 b1out_1 0.18fF
C1000 4bitadder_0/XOR_3/out a3out_0 2.19fF
C1001 4bitadder_0/fulladder_3/and_1/w_26_9# 4bitadder_0/fulladder_3/or_0/b 0.03fF
C1002 comparator_0/not_6/w_n2_10# comparator_0/a2bar 0.03fF
C1003 4bitadder_0/fulladder_1/and_0/w_26_9# vdd 0.03fF
C1004 vdd 4bitadder_1/fulladder_1/axorb 0.15fF
C1005 b2out_2 comparator_0/xnor_1/XOR_0/bbar 0.02fF
C1006 4bitadder_0/fulladder_2/XOR_0/w_62_37# a2out_0 0.02fF
C1007 b0 vdd 0.47fF
C1008 AND_Block_0/and_1/w_n43_8# b1out_3 0.09fF
C1009 4bitadder_0/fulladder_2/axorb 4bitadder_0/fulladder_2/and_0/w_n43_8# 0.09fF
C1010 4bitadder_0/fulladder_2/or_0/w_n48_101# vdd 0.05fF
C1011 vdd comparator_0/not_6/w_n2_10# 0.18fF
C1012 4bitadder_0/fulladder_0/or_0/w_58_101# 4bitadder_0/c1 0.02fF
C1013 a3 b0 0.37fF
C1014 4bitadder_0/fulladder_2/XOR_0/bbar 4bitadder_0/XOR_2/out 0.02fF
C1015 a1out_2 boout_2 0.64fF
C1016 b1out_2 a0out_2 1.11fF
C1017 a0out_3 vdd 0.13fF
C1018 4bitadder_0/XOR_2/out 4bitadder_0/XOR_2/w_62_n20# 0.04fF
C1019 comparator_0/5input_AND_0/not_0/in comparator_0/5input_AND_0/w_106_n113# 0.03fF
C1020 enable_0/and_7/w_n43_8# enable_0/en 0.09fF
C1021 vdd 4bitadder_1/fulladder_1/and_1/w_n43_8# 0.07fF
C1022 enable_3/en enable_3/and_6/w_n43_8# 0.09fF
C1023 4bitadder_1/XOR_1/w_62_n20# 4bitadder_1/XOR_1/bbar 0.13fF
C1024 4bitadder_1/b0xorM 4bitadder_1/XOR_0/w_62_37# 0.02fF
C1025 comparator_0/5input_AND_1/not_0/in gnd 0.10fF
C1026 comparator_0/5input_AND_0/not_0/in comparator_0/a3xnorb3 0.23fF
C1027 a3out_2 gnd 0.76fF
C1028 4bitadder_1/fulladder_3/XOR_1/w_62_37# s3_sub 0.02fF
C1029 comparator_0/xnor_0/XOR_0/w_62_37# b3out_2 0.13fF
C1030 4bitadder_1/fulladder_2/XOR_0/w_62_n20# 4bitadder_1/fulladder_2/XOR_0/abar 0.02fF
C1031 4bitadder_0/fulladder_2/XOR_1/w_16_n1# 4bitadder_0/fulladder_2/XOR_1/bbar 0.03fF
C1032 4bitadder_0/fulladder_2/XOR_1/w_62_n20# s2_add 0.04fF
C1033 4bitadder_0/fulladder_2/XOR_1/w_n34_n1# 4bitadder_0/fulladder_2/XOR_1/abar 0.03fF
C1034 4bitadder_0/fulladder_0/and_0/a_n26_14# s0 0.10fF
C1035 enable_2/and_6/w_26_9# b2out_2 0.03fF
C1036 4bitadder_1/XOR_3/out 4bitadder_1/XOR_3/w_62_n20# 0.04fF
C1037 4bitadder_0/fulladder_0/axorb vdd 0.15fF
C1038 gnd 4bitadder_1/XOR_2/abar 0.13fF
C1039 4bitadder_1/fulladder_1/XOR_0/w_62_37# a1out_1 0.02fF
C1040 b3out_2 comparator_0/xnor_0/not_0/in 0.13fF
C1041 a3out_2 comparator_0/xnor_0/XOR_0/abar 0.13fF
C1042 vdd comparator_0/5input_AND_0/w_n37_15# 0.05fF
C1043 gnd 4bitadder_1/XOR_0/abar 0.15fF
C1044 vdd 4bitadder_1/fulladder_2/XOR_0/w_16_n1# 0.02fF
C1045 enable_3/and_0/w_n43_8# enable_3/and_0/a_n26_14# 0.02fF
C1046 4bitadder_1/fulladder_1/XOR_0/w_62_n20# 4bitadder_1/fulladder_1/XOR_0/abar 0.02fF
C1047 4bitadder_0/fulladder_2/XOR_1/w_n34_n1# vdd 0.02fF
C1048 enable_2/and_3/w_26_9# a3out_2 0.03fF
C1049 comparator_0/5input_AND_1/not_0/in comparator_0/5input_AND_1/not_0/w_n2_10# 0.09fF
C1050 vdd b3out_2 0.82fF
C1051 vdd comparator_0/t4 0.04fF
C1052 comparator_0/4input_AND_0/not_0/w_n2_10# equal 0.03fF
C1053 a1out_1 a2out_1 7.75fF
C1054 vdd b2out_1 0.05fF
C1055 vdd 4bitadder_1/XOR_1/w_16_n1# 0.02fF
C1056 comparator_0/b3bar gnd 0.27fF
C1057 enable_0/and_1/w_n43_8# enable_0/and_1/a_n26_14# 0.02fF
C1058 comparator_0/a1xnorb1 comparator_0/5input_AND_0/not_0/in 0.23fF
C1059 AND_Block_0/and_3/w_n43_8# vdd 0.07fF
C1060 comparator_0/4input_AND_0/not_0/in comparator_0/4input_AND_0/w_68_n95# 0.02fF
C1061 comparator_0/xnor_2/XOR_0/abar gnd 0.14fF
C1062 4bitadder_0/fulladder_3/and_0/w_n43_8# vdd 0.07fF
C1063 4bitadder_0/b0xorM a0out_0 1.79fF
C1064 4bitadder_0/fulladder_0/and_1/w_26_9# 4bitadder_0/fulladder_0/or_0/b 0.03fF
C1065 enable_0/and_5/w_26_9# enable_0/and_5/a_n26_14# 0.09fF
C1066 enable_2/and_7/a_n26_14# b3 0.31fF
C1067 b2out_0 4bitadder_0/XOR_1/abar 1.51fF
C1068 enable_3/and_3/w_26_9# a3out_3 0.03fF
C1069 comparator_0/a1xnorb1 comparator_0/5input_AND_0/w_106_n113# 0.17fF
C1070 4bitadder_0/c1 4bitadder_0/fulladder_1/XOR_1/w_62_37# 0.13fF
C1071 enable_0/en b2 0.38fF
C1072 b2out_0 gnd 1.03fF
C1073 a3out_2 comparator_0/a2xnorb2 0.15fF
C1074 comparator_0/5input_AND_1/not_0/in comparator_0/a2xnorb2 0.23fF
C1075 a2out_2 a0out_2 0.55fF
C1076 vdd comparator_0/t3 0.04fF
C1077 comparator_0/a1xnorb1 comparator_0/a3xnorb3 1.11fF
C1078 4bitadder_0/XOR_1/w_62_n20# 4bitadder_0/XOR_1/bbar 0.13fF
C1079 enable_2/and_3/a_n26_14# a3 0.31fF
C1080 enable_1/and_7/w_26_9# enable_1/and_7/a_n26_14# 0.09fF
C1081 vdd a1out_2 1.25fF
C1082 comparator_0/not_3/w_n2_10# comparator_0/b3bar 0.03fF
C1083 4bitadder_0/fulladder_3/XOR_1/w_62_37# s3_add 0.02fF
C1084 4bitadder_0/c1 s1_add 0.04fF
C1085 4bitadder_0/fulladder_0/or_0/w_n48_101# vdd 0.05fF
C1086 4bitadder_0/fulladder_3/XOR_0/abar gnd 0.15fF
C1087 4bitadder_0/fulladder_2/XOR_0/w_62_n20# 4bitadder_0/fulladder_2/XOR_0/abar 0.02fF
C1088 comparator_0/a0bar comparator_0/a2xnorb2 0.41fF
C1089 4bitadder_1/fulladder_2/axorb 4bitadder_1/fulladder_2/XOR_1/abar 0.13fF
C1090 4bitadder_0/XOR_3/out s0 0.16fF
C1091 enable_1/and_7/w_26_9# b3out_1 0.03fF
C1092 enable_0/and_6/w_26_9# vdd 0.03fF
C1093 comparator_0/4input_AND_2/not_0/in comparator_0/4input_AND_2/w_n47_52# 0.02fF
C1094 4bitadder_0/XOR_3/out 4bitadder_0/XOR_3/w_62_n20# 0.04fF
C1095 decoder_0/and_3/w_n43_8# s1 0.09fF
C1096 4bitadder_0/fulladder_0/and_0/w_n43_8# vdd 0.07fF
C1097 enable_0/and_7/w_n43_8# b3 0.09fF
C1098 b1out_2 comparator_0/4input_AND_2/not_0/in 0.18fF
C1099 vdd comparator_0/xnor_3/XOR_0/w_n34_n1# 0.02fF
C1100 4bitadder_1/fulladder_2/and_0/a_n26_14# 4bitadder_1/fulladder_2/and_0/w_n43_8# 0.02fF
C1101 vdd 4bitadder_1/fulladder_0/and_1/w_n43_8# 0.07fF
C1102 gnd 4bitadder_1/fulladder_2/or_0/a 0.01fF
C1103 4bitadder_0/fulladder_0/axorb s0 0.54fF
C1104 enable_0/and_4/w_26_9# b0out_0 0.03fF
C1105 4bitadder_1/fulladder_3/or_0/a_n15_32# 4bitadder_1/fulladder_3/or_0/b 0.19fF
C1106 comparator_0/b3bar comparator_0/a2xnorb2 0.12fF
C1107 comparator_0/t5 comparator_0/t6 0.21fF
C1108 vdd comparator_0/a0xnorb0 0.04fF
C1109 4bitadder_1/fulladder_1/axorb 4bitadder_1/fulladder_1/and_0/w_n43_8# 0.09fF
C1110 enable_0/en enable_0/and_0/w_n43_8# 0.09fF
C1111 b0out_0 4bitadder_0/XOR_0/abar 0.13fF
C1112 s0 b2out_1 0.35fF
C1113 4bitadder_0/fulladder_2/and_1/w_n43_8# vdd 0.07fF
C1114 4bitadder_0/fulladder_1/and_1/w_n43_8# a1out_0 0.09fF
C1115 comparator_0/a1bar comparator_0/4input_AND_2/w_n47_52# 0.16fF
C1116 enable_1/and_1/w_n43_8# a1 0.09fF
C1117 4bitadder_1/XOR_1/w_16_n1# s0 0.11fF
C1118 4bitadder_1/fulladder_0/and_0/a_n26_14# s0 0.10fF
C1119 comparator_0/a1bar b1out_2 0.44fF
C1120 comparator_0/3input_AND_0/not_0/in comparator_0/3input_AND_0/not_0/w_n2_10# 0.09fF
C1121 comparator_0/xnor_2/not_0/w_n2_10# comparator_0/xnor_2/not_0/in 0.09fF
C1122 4bitadder_0/fulladder_1/or_0/a vdd 0.14fF
C1123 4bitadder_0/fulladder_0/XOR_0/abar gnd 0.15fF
C1124 comparator_0/4input_OR_0/y gnd 0.03fF
C1125 gnd a1out_1 0.92fF
C1126 4bitadder_1/fulladder_2/or_0/a_n15_32# 4bitadder_1/fulladder_2/or_0/w_n48_101# 0.05fF
C1127 4bitadder_0/b0xorM s0 0.26fF
C1128 4bitadder_0/c2 gnd 0.97fF
C1129 gnd 4bitadder_1/fulladder_3/axorb 0.09fF
C1130 comparator_0/xnor_1/not_0/in gnd 0.03fF
C1131 4bitadder_0/XOR_3/w_16_n1# vdd 0.02fF
C1132 b2 a1 0.31fF
C1133 comparator_0/5input_AND_1/not_0/in comparator_0/5input_AND_1/w_n37_15# 0.05fF
C1134 enable_3/and_1/w_n43_8# enable_3/and_1/a_n26_14# 0.02fF
C1135 4bitadder_1/XOR_3/w_n34_n1# b3out_1 0.11fF
C1136 4bitadder_1/c3 4bitadder_1/fulladder_3/XOR_1/bbar 0.02fF
C1137 4bitadder_0/fulladder_2/and_0/a_n26_14# 4bitadder_0/c2 0.10fF
C1138 b2out_2 comparator_0/a3xnorb3 0.19fF
C1139 4bitadder_0/fulladder_2/axorb 4bitadder_0/fulladder_2/XOR_1/abar 0.13fF
C1140 comparator_0/a0bar comparator_0/5input_AND_1/w_n37_15# 0.17fF
C1141 vdd s2_sub 0.19fF
C1142 vdd comparator_0/xnor_1/XOR_0/w_16_n1# 0.02fF
C1143 b2 b3 0.33fF
C1144 4bitadder_1/XOR_3/w_62_n20# 4bitadder_1/XOR_3/abar 0.02fF
C1145 4bitadder_1/c2 4bitadder_1/XOR_2/out 0.55fF
C1146 enable_0/and_2/w_n43_8# enable_0/and_2/a_n26_14# 0.02fF
C1147 vdd 4bitadder_1/fulladder_1/and_1/w_26_9# 0.03fF
C1148 4bitadder_0/fulladder_2/axorb vdd 0.15fF
C1149 4bitadder_0/fulladder_0/and_0/w_n43_8# s0 0.09fF
C1150 4bitadder_1/fulladder_1/and_1/w_26_9# 4bitadder_1/fulladder_1/or_0/b 0.03fF
C1151 vdd comparator_0/5input_AND_1/w_106_n113# 0.04fF
C1152 enable_2/and_5/w_26_9# vdd 0.03fF
C1153 4bitadder_0/fulladder_0/XOR_1/w_62_37# s0_add 0.02fF
C1154 4bitadder_0/fulladder_3/or_0/a_n15_32# 4bitadder_0/fulladder_3/or_0/b 0.19fF
C1155 enable_0/and_7/w_n43_8# vdd 0.07fF
C1156 b1out_1 b2out_1 0.26fF
C1157 4bitadder_1/fulladder_1/XOR_1/w_62_n20# 4bitadder_1/fulladder_1/XOR_1/bbar 0.13fF
C1158 4bitadder_1/fulladder_0/XOR_0/abar 4bitadder_1/fulladder_0/XOR_0/w_n34_n1# 0.03fF
C1159 comparator_0/3input_AND_1/not_0/in gnd 0.21fF
C1160 vdd comparator_0/not_4/w_n2_10# 0.26fF
C1161 enable_1/and_5/a_n26_14# b1 0.31fF
C1162 a2out_2 comparator_0/3input_AND_0/not_0/in 0.19fF
C1163 comparator_0/4input_OR_0/w_n58_n43# comparator_0/t5 0.13fF
C1164 enable_1/and_7/w_26_9# vdd 0.03fF
C1165 4bitadder_1/fulladder_3/and_1/w_n43_8# 4bitadder_1/fulladder_3/and_1/a_n26_14# 0.02fF
C1166 enable_2/and_4/a_n26_14# b0 0.31fF
C1167 enable_1/and_2/w_26_9# a2out_1 0.03fF
C1168 b2out_2 comparator_0/a1xnorb1 0.27fF
C1169 4bitadder_1/fulladder_0/XOR_1/w_62_37# s0_sub 0.02fF
C1170 decoder_0/and_0/a_n26_14# decoder_0/and_1/b 0.33fF
C1171 comparator_0/3input_AND_0/w_69_n71# comparator_0/a3xnorb3 0.16fF
C1172 vdd comparator_0/4input_AND_0/not_0/w_n2_10# 0.18fF
C1173 comparator_0/4input_AND_1/not_0/in comparator_0/4input_AND_1/w_68_n95# 0.02fF
C1174 enable_0/and_1/w_26_9# vdd 0.03fF
C1175 4bitadder_1/c2 4bitadder_1/fulladder_2/and_0/w_n43_8# 0.09fF
C1176 4bitadder_1/XOR_1/out 4bitadder_1/XOR_1/w_62_37# 0.02fF
C1177 vdd comparator_0/4input_AND_0/w_29_n46# 0.02fF
C1178 4bitadder_0/fulladder_2/XOR_0/w_n34_n1# vdd 0.02fF
C1179 4bitadder_0/fulladder_1/XOR_0/w_n34_n1# a1out_0 0.11fF
C1180 4bitadder_0/fulladder_1/XOR_0/w_16_n1# 4bitadder_0/XOR_1/out 0.11fF
C1181 4bitadder_1/fulladder_0/or_0/a_n15_32# 4bitadder_1/fulladder_0/or_0/w_58_101# 0.13fF
C1182 4bitadder_0/XOR_3/w_16_n1# s0 0.11fF
C1183 4bitadder_0/c3 4bitadder_0/fulladder_3/XOR_1/bbar 0.02fF
C1184 4bitadder_0/fulladder_3/XOR_1/w_16_n1# vdd 0.02fF
C1185 gnd a2out_1 1.13fF
C1186 comparator_0/and_1/a_n26_14# gnd 0.02fF
C1187 vdd comparator_0/t2 0.04fF
C1188 enable_1/en gnd 0.13fF
C1189 4bitadder_0/fulladder_1/XOR_0/abar 4bitadder_0/XOR_1/out 0.25fF
C1190 AND_Block_0/and_0/w_n43_8# a0out_3 0.09fF
C1191 a0_out1 4bitadder_1/b0xorM 1.79fF
C1192 4bitadder_0/XOR_3/abar s0 0.30fF
C1193 enable_1/and_1/w_n43_8# vdd 0.07fF
C1194 enable_0/en enable_0/and_2/w_n43_8# 0.09fF
C1195 4bitadder_0/c2 4bitadder_0/XOR_2/out 0.55fF
C1196 4bitadder_0/XOR_3/w_62_n20# 4bitadder_0/XOR_3/abar 0.02fF
C1197 comparator_0/3input_AND_0/not_0/in comparator_0/3input_AND_0/w_n14_24# 0.03fF
C1198 a0out_2 comparator_0/5input_AND_0/w_n37_15# 0.17fF
C1199 a0out_3 b0out_3 2.02fF
C1200 enable_3/and_5/a_n26_14# enable_3/and_5/w_26_9# 0.09fF
C1201 enable_1/and_6/w_n43_8# vdd 0.07fF
C1202 b2 vdd 0.45fF
C1203 4bitadder_0/XOR_0/w_n34_n1# vdd 0.02fF
C1204 a1out_0 vdd 0.28fF
C1205 fc_sub 4bitadder_1/fulladder_3/or_0/w_58_101# 0.02fF
C1206 gnd 4bitadder_1/fulladder_1/XOR_1/abar 0.15fF
C1207 vdd 4bitadder_1/XOR_3/w_n34_n1# 0.02fF
C1208 b3out_2 a0out_2 0.58fF
C1209 a3out_2 boout_2 0.37fF
C1210 boout_2 comparator_0/5input_AND_1/not_0/in 0.23fF
C1211 4bitadder_0/fulladder_1/XOR_1/w_62_n20# 4bitadder_0/fulladder_1/XOR_1/bbar 0.13fF
C1212 enable_3/and_1/w_26_9# vdd 0.03fF
C1213 enable_3/and_7/w_26_9# b3out_3 0.03fF
C1214 comparator_0/and_1/w_n43_8# comparator_0/and_1/a_n26_14# 0.02fF
C1215 comparator_0/and_1/w_26_9# comparator_0/t1 0.03fF
C1216 enable_1/and_6/w_26_9# vdd 0.03fF
C1217 b2 a3 0.31fF
C1218 comparator_0/xnor_1/XOR_0/w_n34_n1# a2out_2 0.11fF
C1219 enable_3/en enable_3/and_1/w_n43_8# 0.09fF
C1220 b1out_3 gnd 0.25fF
C1221 4bitadder_1/fulladder_1/XOR_0/bbar 4bitadder_1/fulladder_1/XOR_0/w_16_n1# 0.03fF
C1222 4bitadder_0/fulladder_3/and_1/w_n43_8# 4bitadder_0/fulladder_3/and_1/a_n26_14# 0.02fF
C1223 4bitadder_0/fulladder_2/or_0/w_n48_101# 4bitadder_0/fulladder_2/or_0/a_n15_32# 0.05fF
C1224 enable_2/and_5/a_n26_14# enable_2/and_5/w_26_9# 0.09fF
C1225 enable_3/and_2/w_n43_8# enable_3/and_2/a_n26_14# 0.02fF
C1226 comparator_0/a0xnorb0 comparator_0/4input_AND_0/w_68_n95# 0.16fF
C1227 comparator_0/a0bar boout_2 0.33fF
C1228 4bitadder_0/fulladder_0/XOR_1/w_16_n1# vdd 0.02fF
C1229 vdd 4bitadder_1/fulladder_2/and_0/w_26_9# 0.03fF
C1230 enable_0/and_3/w_26_9# a3out_0 0.03fF
C1231 4bitadder_1/c3 4bitadder_1/fulladder_3/axorb 0.60fF
C1232 comparator_0/xnor_1/XOR_0/w_62_n20# comparator_0/xnor_1/XOR_0/abar 0.02fF
C1233 4bitadder_1/fulladder_0/and_1/a_n26_14# 4bitadder_1/fulladder_0/and_1/w_26_9# 0.09fF
C1234 enable_1/and_1/w_n43_8# enable_1/and_1/a_n26_14# 0.02fF
C1235 enable_3/and_0/w_26_9# a0out_3 0.03fF
C1236 4bitadder_0/c2 4bitadder_0/fulladder_2/and_0/w_n43_8# 0.09fF
C1237 comparator_0/5input_AND_0/not_0/w_n2_10# comparator_0/5input_AND_0/not_0/in 0.09fF
C1238 enable_0/and_3/w_n43_8# enable_0/and_3/a_n26_14# 0.02fF
C1239 b1out_3 a3out_3 0.11fF
C1240 vdd 4bitadder_1/fulladder_3/or_0/w_n48_101# 0.05fF
C1241 vdd 4bitadder_1/fulladder_0/XOR_1/w_n34_n1# 0.02fF
C1242 b1 a0 0.28fF
C1243 decoder_0/and_1/b decoder_0/not_1/w_n2_10# 0.03fF
C1244 a1out_2 a0out_2 0.58fF
C1245 4bitadder_0/fulladder_3/or_0/b gnd 0.37fF
C1246 4bitadder_1/fulladder_0/XOR_1/w_n34_n1# 4bitadder_1/fulladder_0/axorb 0.11fF
C1247 enable_3/en enable_3/and_5/w_n43_8# 0.09fF
C1248 comparator_0/5input_AND_0/not_0/in comparator_0/5input_AND_0/w_31_n55# 0.03fF
C1249 4bitadder_0/fulladder_1/or_0/w_58_101# vdd 0.05fF
C1250 enable_0/and_0/w_n43_8# vdd 0.07fF
C1251 4bitadder_1/fulladder_3/XOR_0/abar a3out_1 0.13fF
C1252 4bitadder_0/XOR_1/abar gnd 0.23fF
C1253 comparator_0/b1bar comparator_0/4input_AND_1/w_n8_2# 0.16fF
C1254 comparator_0/xnor_3/XOR_0/w_n34_n1# a0out_2 0.11fF
C1255 b0out_0 a2out_0 0.12fF
C1256 enable_3/en b1 0.25fF
C1257 comparator_0/b1bar comparator_0/a3xnorb3 0.35fF
C1258 4bitadder_0/fulladder_3/and_1/w_26_9# vdd 0.03fF
C1259 4bitadder_1/fulladder_2/XOR_0/w_16_n1# 4bitadder_1/fulladder_2/XOR_0/bbar 0.03fF
C1260 4bitadder_1/fulladder_2/XOR_0/w_n34_n1# 4bitadder_1/fulladder_2/XOR_0/abar 0.03fF
C1261 comparator_0/xnor_0/XOR_0/w_62_37# a3out_2 0.02fF
C1262 enable_2/en decoder_0/and_2/w_26_9# 0.03fF
C1263 4bitadder_1/fulladder_0/XOR_0/w_62_n20# 4bitadder_1/fulladder_0/XOR_0/abar 0.02fF
C1264 fc_add 4bitadder_0/fulladder_3/or_0/w_58_101# 0.02fF
C1265 a2out_2 comparator_0/b2bar 0.44fF
C1266 comparator_0/5input_AND_0/w_31_n55# comparator_0/a3xnorb3 0.21fF
C1267 comparator_0/xnor_0/XOR_0/abar gnd 0.14fF
C1268 AND_Block_0/and_2/w_26_9# vdd 0.03fF
C1269 enable_0/and_3/w_26_9# vdd 0.03fF
C1270 a1out_0 s0 2.21fF
C1271 4bitadder_1/fulladder_3/XOR_1/w_62_n20# 4bitadder_1/fulladder_3/XOR_1/abar 0.02fF
C1272 4bitadder_1/fulladder_0/XOR_1/w_62_n20# 4bitadder_1/fulladder_0/XOR_1/abar 0.02fF
C1273 comparator_0/xnor_0/XOR_0/w_62_n20# comparator_0/xnor_0/XOR_0/bbar 0.13fF
C1274 vdd comparator_0/t8 0.04fF
C1275 a3out_3 gnd 0.14fF
C1276 vdd 4bitadder_1/fulladder_3/XOR_1/w_n34_n1# 0.02fF
C1277 vdd comparator_0/3input_AND_1/w_32_n21# 0.03fF
C1278 4bitadder_0/fulladder_0/or_0/b gnd 0.37fF
C1279 vdd a3out_2 0.91fF
C1280 s0 4bitadder_1/XOR_3/bbar 0.02fF
C1281 vdd 4bitadder_1/XOR_2/w_16_n1# 0.02fF
C1282 4bitadder_0/c3 4bitadder_0/fulladder_3/axorb 0.60fF
C1283 4bitadder_0/fulladder_0/XOR_1/w_16_n1# s0 0.11fF
C1284 enable_3/and_0/w_n43_8# vdd 0.07fF
C1285 vdd comparator_0/4input_AND_1/w_29_n46# 0.02fF
C1286 enable_0/en enable_0/and_4/w_n43_8# 0.09fF
C1287 b2out_0 a3out_0 0.11fF
C1288 b0out_1 4bitadder_1/XOR_0/abar 0.13fF
C1289 vdd 4bitadder_1/fulladder_1/or_0/w_58_101# 0.05fF
C1290 4bitadder_1/XOR_1/out 4bitadder_1/c1 0.37fF
C1291 vdd comparator_0/a0bar 0.30fF
C1292 AND_Block_0/and_3/w_26_9# AND_Block_0/and_3/a_n26_14# 0.09fF
C1293 comparator_0/t8 comparator_0/t6 0.29fF
C1294 comparator_0/4input_AND_0/not_0/in comparator_0/4input_AND_0/w_n8_2# 0.02fF
C1295 comparator_0/xnor_2/not_0/in gnd 0.03fF
C1296 comparator_0/b1bar comparator_0/not_1/w_n2_10# 0.03fF
C1297 4bitadder_0/fulladder_2/or_0/w_n48_101# 4bitadder_0/fulladder_2/or_0/b 0.12fF
C1298 4bitadder_0/fulladder_0/XOR_1/abar s0 0.27fF
C1299 4bitadder_0/fulladder_0/and_1/w_n43_8# 4bitadder_0/fulladder_0/and_1/a_n26_14# 0.02fF
C1300 4bitadder_0/fulladder_0/and_1/w_26_9# vdd 0.03fF
C1301 AND_Block_0/and_1/w_n43_8# vdd 0.07fF
C1302 a1out_1 b3out_1 0.24fF
C1303 4bitadder_1/fulladder_1/and_0/a_n26_14# 4bitadder_1/fulladder_1/and_0/w_26_9# 0.09fF
C1304 comparator_0/a2xnorb2 gnd 1.27fF
C1305 comparator_0/4input_AND_2/w_n47_52# comparator_0/a3xnorb3 0.04fF
C1306 comparator_0/3input_AND_0/w_n14_24# comparator_0/b2bar 0.16fF
C1307 4bitadder_0/fulladder_3/XOR_0/abar a3out_0 0.13fF
C1308 comparator_0/5input_AND_0/w_68_n82# comparator_0/a2xnorb2 0.16fF
C1309 enable_3/and_3/w_26_9# vdd 0.03fF
C1310 4bitadder_1/fulladder_2/axorb 4bitadder_1/fulladder_2/XOR_1/w_62_37# 0.02fF
C1311 4bitadder_1/c2 4bitadder_1/fulladder_2/XOR_1/w_16_n1# 0.11fF
C1312 b1out_2 comparator_0/a3xnorb3 0.36fF
C1313 4bitadder_0/fulladder_1/and_0/a_n26_14# 4bitadder_0/fulladder_1/and_0/w_26_9# 0.09fF
C1314 enable_3/en enable_3/and_3/w_n43_8# 0.09fF
C1315 vdd comparator_0/xnor_2/XOR_0/w_16_n1# 0.02fF
C1316 vdd comparator_0/b3bar 0.04fF
C1317 4bitadder_0/fulladder_2/XOR_0/w_16_n1# 4bitadder_0/fulladder_2/XOR_0/bbar 0.03fF
C1318 4bitadder_0/fulladder_2/XOR_0/w_n34_n1# 4bitadder_0/fulladder_2/XOR_0/abar 0.03fF
C1319 enable_3/and_3/w_n43_8# enable_3/and_3/a_n26_14# 0.02fF
C1320 4bitadder_1/c2 4bitadder_1/fulladder_2/XOR_1/abar 0.27fF
C1321 vdd comparator_0/4input_AND_2/w_68_n95# 0.02fF
C1322 enable_2/en b1 0.30fF
C1323 4bitadder_1/fulladder_0/XOR_1/w_62_n20# 4bitadder_1/fulladder_0/XOR_1/bbar 0.13fF
C1324 4bitadder_0/fulladder_3/XOR_1/w_62_n20# 4bitadder_0/fulladder_3/XOR_1/abar 0.02fF
C1325 comparator_0/xnor_2/XOR_0/w_62_37# comparator_0/xnor_2/not_0/in 0.02fF
C1326 comparator_0/not_4/w_n2_10# a0out_2 0.09fF
C1327 4bitadder_1/fulladder_2/or_0/w_58_101# 4bitadder_1/c3 0.02fF
C1328 b2out_0 vdd 0.05fF
C1329 4bitadder_0/fulladder_3/XOR_0/w_16_n1# vdd 0.02fF
C1330 4bitadder_0/XOR_2/out gnd 0.42fF
C1331 enable_0/and_4/w_n43_8# enable_0/and_4/a_n26_14# 0.02fF
C1332 vdd 4bitadder_1/fulladder_0/and_0/w_26_9# 0.03fF
C1333 b1 a2 0.28fF
C1334 s1 decoder_0/and_3/a_n26_14# 0.31fF
C1335 enable_0/and_7/a_n26_14# b3 0.31fF
C1336 vdd comparator_0/xnor_3/not_0/w_n2_10# 0.18fF
C1337 enable_1/en enable_1/and_3/w_n43_8# 0.09fF
C1338 gnd decoder_0/and_1/b 0.19fF
C1339 4bitadder_1/fulladder_3/and_0/w_26_9# 4bitadder_1/fulladder_3/or_0/a 0.03fF
C1340 4bitadder_1/fulladder_0/or_0/w_n48_101# 4bitadder_1/fulladder_0/or_0/a 0.12fF
C1341 vdd comparator_0/xnor_2/not_0/w_n2_10# 0.18fF
C1342 comparator_0/4input_OR_0/NOT_0/w_n2_10# agb 0.03fF
C1343 b1out_2 comparator_0/xnor_2/XOR_0/bbar 0.02fF
C1344 4bitadder_0/fulladder_0/axorb 4bitadder_0/fulladder_0/XOR_0/w_62_n20# 0.04fF
C1345 enable_1/and_6/a_n26_14# enable_1/and_6/w_n43_8# 0.02fF
C1346 enable_0/and_2/w_n43_8# vdd 0.07fF
C1347 comparator_0/a1xnorb1 b1out_2 0.69fF
C1348 4bitadder_1/fulladder_1/or_0/w_58_101# 4bitadder_1/fulladder_1/or_0/a_n15_32# 0.13fF
C1349 enable_2/and_0/w_n43_8# a0 0.09fF
C1350 enable_1/and_6/a_n26_14# b2 0.31fF
C1351 s0 4bitadder_1/XOR_2/w_16_n1# 0.11fF
C1352 comparator_0/not_1/w_n2_10# b1out_2 0.09fF
C1353 vdd 4bitadder_1/fulladder_3/and_1/w_n43_8# 0.07fF
C1354 enable_1/and_6/a_n26_14# enable_1/and_6/w_26_9# 0.09fF
C1355 4bitadder_1/fulladder_2/and_1/w_26_9# 4bitadder_1/fulladder_2/and_1/a_n26_14# 0.09fF
C1356 4bitadder_1/fulladder_1/XOR_0/bbar 4bitadder_1/XOR_1/out 0.02fF
C1357 comparator_0/b0bar comparator_0/a2xnorb2 0.38fF
C1358 vdd 4bitadder_1/fulladder_2/or_0/a 0.14fF
C1359 comparator_0/4input_OR_0/w_n58_n43# comparator_0/t8 0.13fF
C1360 s0 4bitadder_1/XOR_2/abar 0.28fF
C1361 a1out_0 4bitadder_0/fulladder_1/and_1/a_n26_14# 0.10fF
C1362 4bitadder_1/XOR_1/w_n34_n1# 4bitadder_1/XOR_1/abar 0.03fF
C1363 4bitadder_1/XOR_0/abar s0 1.07fF
C1364 gnd 4bitadder_1/c3 0.91fF
C1365 4bitadder_0/fulladder_2/axorb 4bitadder_0/fulladder_2/XOR_1/w_62_37# 0.02fF
C1366 4bitadder_0/c2 4bitadder_0/fulladder_2/XOR_1/w_16_n1# 0.11fF
C1367 b1 enable_0/and_5/w_n43_8# 0.09fF
C1368 a2out_1 b3out_1 0.33fF
C1369 enable_2/and_5/w_n43_8# vdd 0.07fF
C1370 4bitadder_0/fulladder_0/XOR_0/w_16_n1# vdd 0.02fF
C1371 enable_1/en a1 0.28fF
C1372 a2out_2 comparator_0/a3xnorb3 0.60fF
C1373 comparator_0/4input_OR_0/NOT_0/w_n2_10# vdd 0.18fF
C1374 4bitadder_0/c2 4bitadder_0/fulladder_2/XOR_1/abar 0.27fF
C1375 a1out_1 b0out_1 0.11fF
C1376 enable_0/en gnd 0.01fF
C1377 4bitadder_1/fulladder_3/or_0/a_n15_32# 4bitadder_1/fulladder_3/or_0/w_58_101# 0.13fF
C1378 4bitadder_1/fulladder_1/XOR_0/abar a1out_1 0.13fF
C1379 enable_3/and_2/w_n43_8# vdd 0.07fF
C1380 4bitadder_1/XOR_3/w_16_n1# 4bitadder_1/XOR_3/bbar 0.03fF
C1381 4bitadder_1/XOR_3/w_n34_n1# 4bitadder_1/XOR_3/abar 0.03fF
C1382 4bitadder_0/fulladder_2/and_0/a_n26_14# 4bitadder_0/fulladder_2/and_0/w_n43_8# 0.02fF
C1383 4bitadder_0/fulladder_0/XOR_0/abar a0out_0 0.13fF
C1384 vdd a1out_1 0.33fF
C1385 4bitadder_0/c2 vdd 0.17fF
C1386 4bitadder_0/c1 a1out_0 0.35fF
C1387 4bitadder_0/fulladder_2/or_0/w_58_101# 4bitadder_0/c3 0.02fF
C1388 4bitadder_0/fulladder_1/or_0/w_n48_101# 4bitadder_0/fulladder_1/or_0/a_n15_32# 0.05fF
C1389 enable_1/en b3 0.21fF
C1390 vdd 4bitadder_1/fulladder_3/axorb 0.15fF
C1391 vdd comparator_0/5input_AND_1/w_31_n55# 0.06fF
C1392 4bitadder_0/fulladder_3/or_0/a gnd 0.01fF
C1393 b2out_0 s0 0.30fF
C1394 4bitadder_0/fulladder_3/and_0/w_26_9# 4bitadder_0/fulladder_3/or_0/a 0.03fF
C1395 enable_2/and_7/w_n43_8# b3 0.09fF
C1396 4bitadder_0/fulladder_0/XOR_1/w_62_n20# 4bitadder_0/fulladder_0/XOR_1/abar 0.02fF
C1397 4bitadder_0/fulladder_0/and_0/w_26_9# 4bitadder_0/fulladder_0/and_0/a_n26_14# 0.09fF
C1398 b2 enable_3/and_6/w_n43_8# 0.09fF
C1399 4bitadder_1/fulladder_3/and_1/w_n43_8# 4bitadder_1/XOR_3/out 0.09fF
C1400 b2out_2 b1out_2 0.42fF
C1401 enable_1/and_0/w_n43_8# enable_1/en 0.09fF
C1402 4bitadder_1/fulladder_0/or_0/w_n48_101# 4bitadder_1/fulladder_0/or_0/b 0.12fF
C1403 a2out_2 comparator_0/a1xnorb1 0.46fF
C1404 comparator_0/4input_OR_0/y comparator_0/t6 0.18fF
C1405 boout_2 comparator_0/xnor_3/XOR_0/bbar 0.02fF
C1406 4bitadder_0/fulladder_2/and_1/w_26_9# 4bitadder_0/fulladder_2/and_1/a_n26_14# 0.09fF
C1407 enable_3/and_4/w_n43_8# enable_3/and_4/a_n26_14# 0.02fF
C1408 comparator_0/4input_AND_1/not_0/in comparator_0/4input_AND_1/w_n8_2# 0.02fF
C1409 vdd comparator_0/and_0/w_26_9# 0.03fF
C1410 comparator_0/4input_AND_1/not_0/in comparator_0/a3xnorb3 0.18fF
C1411 4bitadder_0/XOR_1/w_n34_n1# 4bitadder_0/XOR_1/abar 0.03fF
C1412 4bitadder_0/fulladder_1/XOR_0/w_62_37# 4bitadder_0/XOR_1/out 0.13fF
C1413 vdd comparator_0/4input_AND_0/w_n47_52# 0.02fF
C1414 4bitadder_0/XOR_3/w_62_37# s0 0.13fF
C1415 b2out_3 AND_Block_0/and_2/a_n26_14# 0.31fF
C1416 enable_3/and_5/w_n43_8# enable_3/and_5/a_n26_14# 0.02fF
C1417 vdd enable_2/and_7/w_26_9# 0.03fF
C1418 vdd 4bitadder_1/fulladder_3/XOR_0/w_n34_n1# 0.02fF
C1419 vdd decoder_0/not_1/w_n2_10# 0.18fF
C1420 4bitadder_1/XOR_0/w_62_n20# 4bitadder_1/XOR_0/abar 0.02fF
C1421 enable_2/and_0/w_n43_8# enable_2/en 0.09fF
C1422 b1 b0 4.71fF
C1423 4bitadder_0/fulladder_0/or_0/a gnd 0.01fF
C1424 4bitadder_0/fulladder_3/or_0/a_n15_32# 4bitadder_0/fulladder_3/or_0/w_58_101# 0.13fF
C1425 4bitadder_0/XOR_2/w_n34_n1# vdd 0.02fF
C1426 4bitadder_0/fulladder_0/axorb 4bitadder_0/fulladder_0/XOR_1/w_n34_n1# 0.11fF
C1427 enable_3/and_5/a_n26_14# b1 0.31fF
C1428 enable_0/and_4/w_n43_8# vdd 0.07fF
C1429 4bitadder_0/XOR_3/w_16_n1# 4bitadder_0/XOR_3/bbar 0.03fF
C1430 4bitadder_0/XOR_3/w_n34_n1# 4bitadder_0/XOR_3/abar 0.03fF
C1431 a1 gnd 0.27fF
C1432 s3_add vdd 0.10fF
C1433 enable_2/and_5/w_n43_8# enable_2/and_5/a_n26_14# 0.02fF
C1434 gnd b3out_1 0.62fF
C1435 comparator_0/t4 comparator_0/t1 0.18fF
C1436 comparator_0/a1xnorb1 comparator_0/4input_AND_0/not_0/in 0.18fF
C1437 a2out_1 b0out_1 0.09fF
C1438 4bitadder_1/fulladder_3/axorb 4bitadder_1/XOR_3/out 0.13fF
C1439 4bitadder_0/fulladder_2/or_0/w_n48_101# 4bitadder_0/fulladder_2/or_0/a 0.12fF
C1440 vdd comparator_0/4input_AND_1/not_0/w_n2_10# 0.18fF
C1441 4bitadder_1/fulladder_0/and_1/w_n43_8# 4bitadder_1/b0xorM 0.09fF
C1442 a1out_1 s0 0.21fF
C1443 enable_2/and_1/w_26_9# vdd 0.03fF
C1444 vdd a2out_1 0.33fF
C1445 boout_2 gnd 0.90fF
C1446 b3 gnd 0.29fF
C1447 4bitadder_1/fulladder_2/axorb 4bitadder_1/fulladder_2/XOR_0/w_62_37# 0.02fF
C1448 4bitadder_1/fulladder_0/XOR_1/w_n34_n1# 4bitadder_1/fulladder_0/XOR_1/abar 0.03fF
C1449 a3out_2 a0out_2 0.60fF
C1450 enable_2/and_2/w_26_9# a2out_2 0.03fF
C1451 enable_1/en vdd 0.92fF
C1452 4bitadder_0/fulladder_3/and_1/w_n43_8# 4bitadder_0/XOR_3/out 0.09fF
C1453 4bitadder_0/fulladder_1/axorb gnd 0.09fF
C1454 4bitadder_0/fulladder_1/axorb 4bitadder_0/fulladder_1/XOR_0/w_62_n20# 0.04fF
C1455 4bitadder_0/fulladder_1/or_0/w_n48_101# 4bitadder_0/fulladder_1/or_0/b 0.12fF
C1456 enable_3/and_7/w_n43_8# b3 0.09fF
C1457 4bitadder_1/XOR_1/out 4bitadder_1/fulladder_1/axorb 0.13fF
C1458 comparator_0/t1 comparator_0/t3 0.18fF
C1459 enable_1/en a3 0.28fF
C1460 vdd 4bitadder_1/fulladder_1/XOR_1/w_16_n1# 0.02fF
C1461 enable_2/and_7/w_n43_8# vdd 0.07fF
C1462 a2out_2 b2out_2 0.46fF
C1463 comparator_0/xnor_1/XOR_0/w_16_n1# comparator_0/xnor_1/XOR_0/bbar 0.03fF
C1464 comparator_0/xnor_1/XOR_0/w_62_n20# comparator_0/xnor_1/not_0/in 0.04fF
C1465 comparator_0/xnor_1/XOR_0/w_n34_n1# comparator_0/xnor_1/XOR_0/abar 0.03fF
C1466 comparator_0/4input_OR_0/y comparator_0/4input_OR_0/w_n58_n43# 0.02fF
C1467 enable_0/and_6/w_n43_8# b2 0.09fF
C1468 a2out_3 b1out_3 0.12fF
C1469 comparator_0/4input_OR_1/y comparator_0/t1 0.18fF
C1470 enable_3/and_4/w_n43_8# vdd 0.07fF
C1471 4bitadder_1/c1 4bitadder_1/fulladder_1/XOR_1/bbar 0.02fF
C1472 s0_add vdd 0.19fF
C1473 4bitadder_1/fulladder_3/XOR_0/w_62_37# a3out_1 0.02fF
C1474 4bitadder_1/fulladder_2/or_0/w_n48_101# 4bitadder_1/fulladder_2/or_0/b 0.12fF
C1475 b3out_0 4bitadder_0/XOR_3/abar 0.13fF
C1476 4bitadder_1/fulladder_3/axorb 4bitadder_1/fulladder_3/and_0/w_n43_8# 0.09fF
C1477 4bitadder_0/XOR_0/w_62_n20# 4bitadder_0/XOR_0/abar 0.02fF
C1478 enable_1/and_3/w_26_9# a3out_1 0.03fF
C1479 a3out_0 gnd 0.99fF
C1480 b1out_3 vdd 0.12fF
C1481 4bitadder_1/XOR_1/out 4bitadder_1/fulladder_1/and_1/w_n43_8# 0.09fF
C1482 comparator_0/5input_AND_0/not_0/in comparator_0/5input_AND_0/w_n37_15# 0.05fF
C1483 4bitadder_1/fulladder_3/XOR_0/bbar 4bitadder_1/XOR_3/out 0.02fF
C1484 vdd 4bitadder_1/fulladder_2/or_0/w_58_101# 0.05fF
C1485 4bitadder_0/fulladder_3/axorb 4bitadder_0/XOR_3/out 0.13fF
C1486 enable_0/and_7/w_26_9# enable_0/and_7/a_n26_14# 0.09fF
C1487 boout_2 comparator_0/a2xnorb2 0.69fF
C1488 enable_3/and_6/w_26_9# vdd 0.03fF
C1489 enable_1/and_2/w_26_9# vdd 0.03fF
C1490 a1out_3 a0out_3 23.76fF
C1491 a1out_2 comparator_0/not_5/w_n2_10# 0.09fF
C1492 comparator_0/xnor_3/XOR_0/w_n34_n1# comparator_0/xnor_3/XOR_0/abar 0.03fF
C1493 4bitadder_0/fulladder_1/XOR_0/w_62_n20# 4bitadder_0/fulladder_1/XOR_0/bbar 0.13fF
C1494 enable_2/and_6/w_26_9# enable_2/and_6/a_n26_14# 0.09fF
C1495 comparator_0/xnor_0/not_0/in gnd 0.03fF
C1496 4bitadder_0/XOR_2/bbar s0 0.02fF
C1497 4bitadder_1/fulladder_3/XOR_1/w_16_n1# 4bitadder_1/fulladder_3/XOR_1/bbar 0.03fF
C1498 4bitadder_1/fulladder_3/XOR_1/w_62_n20# s3_sub 0.04fF
C1499 4bitadder_1/fulladder_3/XOR_1/w_n34_n1# 4bitadder_1/fulladder_3/XOR_1/abar 0.03fF
C1500 4bitadder_0/fulladder_2/axorb 4bitadder_0/fulladder_2/XOR_0/w_62_37# 0.02fF
C1501 4bitadder_0/fulladder_2/XOR_1/abar gnd 0.15fF
C1502 a2out_3 gnd 0.17fF
C1503 gnd b0out_1 0.14fF
C1504 a2out_1 s0 0.22fF
C1505 enable_1/en decoder_0/and_1/w_26_9# 0.03fF
C1506 4bitadder_1/XOR_2/w_n34_n1# b2out_1 0.11fF
C1507 gnd 4bitadder_1/fulladder_1/XOR_0/abar 0.15fF
C1508 enable_2/en enable_2/and_1/w_n43_8# 0.09fF
C1509 vdd gnd 5.30fF
C1510 a0out_0 gnd 0.46fF
C1511 gnd 4bitadder_1/fulladder_1/or_0/b 0.37fF
C1512 vdd comparator_0/5input_AND_0/w_68_n82# 0.05fF
C1513 vdd comparator_0/xnor_0/XOR_0/w_16_n1# 0.02fF
C1514 4bitadder_0/fulladder_3/and_0/w_26_9# vdd 0.03fF
C1515 4bitadder_1/XOR_2/w_62_n20# 4bitadder_1/XOR_2/abar 0.02fF
C1516 gnd 4bitadder_1/fulladder_0/axorb 0.09fF
C1517 4bitadder_0/fulladder_0/XOR_1/w_62_37# s0 0.13fF
C1518 vdd comparator_0/4input_AND_1/w_n47_52# 0.02fF
C1519 a2out_3 a3out_3 0.39fF
C1520 a3 gnd 0.27fF
C1521 vdd decoder_0/and_2/w_n43_8# 0.07fF
C1522 4bitadder_0/fulladder_3/XOR_0/w_62_37# a3out_0 0.02fF
C1523 enable_3/and_7/w_n43_8# vdd 0.07fF
C1524 AND_Block_0/and_3/w_n43_8# b3out_3 0.09fF
C1525 4bitadder_1/fulladder_0/and_0/a_n26_14# 4bitadder_1/fulladder_0/and_0/w_n43_8# 0.02fF
C1526 4bitadder_0/fulladder_3/axorb 4bitadder_0/fulladder_3/and_0/w_n43_8# 0.09fF
C1527 s0_add s0 0.04fF
C1528 4bitadder_0/fulladder_0/and_1/w_n43_8# 4bitadder_0/b0xorM 0.09fF
C1529 enable_3/and_7/a_n26_14# enable_3/and_7/w_26_9# 0.09fF
C1530 4bitadder_1/XOR_0/abar 4bitadder_1/XOR_0/w_n34_n1# 0.03fF
C1531 enable_3/en a0 0.23fF
C1532 enable_2/and_3/w_26_9# vdd 0.03fF
C1533 4bitadder_0/fulladder_3/XOR_0/bbar 4bitadder_0/XOR_3/out 0.02fF
C1534 vdd comparator_0/5input_AND_1/not_0/w_n2_10# 0.17fF
C1535 vdd comparator_0/not_3/w_n2_10# 0.18fF
C1536 comparator_0/b0bar comparator_0/5input_AND_0/w_n4_n20# 0.18fF
C1537 4bitadder_1/c2 4bitadder_1/fulladder_2/XOR_1/w_62_37# 0.13fF
C1538 a1out_2 comparator_0/a3xnorb3 0.53fF
C1539 vdd comparator_0/and_1/w_n43_8# 0.07fF
C1540 vdd 4bitadder_1/XOR_0/w_16_n1# 0.02fF
C1541 vdd 4bitadder_1/fulladder_0/or_0/w_58_101# 0.05fF
C1542 b3out_2 comparator_0/a1xnorb1 0.42fF
C1543 4bitadder_0/fulladder_1/axorb 4bitadder_0/fulladder_1/XOR_1/w_n34_n1# 0.11fF
C1544 vdd decoder_0/and_3/w_26_9# 0.03fF
C1545 4bitadder_1/fulladder_2/and_0/a_n26_14# 4bitadder_1/fulladder_2/and_0/w_26_9# 0.09fF
C1546 4bitadder_1/c2 s2_sub 0.04fF
C1547 enable_0/en a1 0.35fF
C1548 vdd comparator_0/4input_AND_2/w_n8_2# 0.02fF
C1549 a2out_1 b1out_1 0.12fF
C1550 4bitadder_1/fulladder_3/XOR_0/w_62_n20# 4bitadder_1/fulladder_3/XOR_0/abar 0.02fF
C1551 comparator_0/4input_AND_2/not_0/w_n2_10# comparator_0/t3 0.03fF
C1552 4bitadder_1/fulladder_0/XOR_0/abar 4bitadder_1/b0xorM 0.25fF
C1553 4bitadder_0/fulladder_3/XOR_1/w_16_n1# 4bitadder_0/fulladder_3/XOR_1/bbar 0.03fF
C1554 4bitadder_0/fulladder_3/XOR_1/w_62_n20# s3_add 0.04fF
C1555 4bitadder_0/fulladder_3/XOR_1/w_n34_n1# 4bitadder_0/fulladder_3/XOR_1/abar 0.03fF
C1556 comparator_0/t2 comparator_0/3input_AND_1/not_0/w_n2_10# 0.03fF
C1557 vdd comparator_0/4input_OR_1/w_n58_n43# 0.03fF
C1558 comparator_0/xnor_2/XOR_0/w_n34_n1# a1out_2 0.11fF
C1559 4bitadder_0/fulladder_0/or_0/w_58_101# 4bitadder_0/fulladder_0/or_0/a_n15_32# 0.13fF
C1560 vdd decoder_0/not_0/w_n2_10# 0.18fF
C1561 4bitadder_1/fulladder_0/axorb 4bitadder_1/fulladder_0/XOR_0/w_62_37# 0.02fF
C1562 vdd comparator_0/a2xnorb2 2.46fF
C1563 vdd comparator_0/b0bar 0.14fF
C1564 comparator_0/a0xnorb0 comparator_0/a3xnorb3 0.29fF
C1565 comparator_0/4input_AND_2/not_0/in comparator_0/4input_AND_2/w_68_n95# 0.02fF
C1566 comparator_0/b3bar comparator_0/and_0/a_n26_14# 0.10fF
C1567 gnd 4bitadder_1/XOR_3/out 0.42fF
C1568 4bitadder_1/fulladder_1/and_0/a_n26_14# 4bitadder_1/fulladder_1/and_0/w_n43_8# 0.02fF
C1569 enable_0/en b3 0.10fF
C1570 comparator_0/xnor_2/XOR_0/w_62_n20# comparator_0/xnor_2/XOR_0/abar 0.02fF
C1571 4bitadder_0/XOR_1/abar s0 0.25fF
C1572 comparator_0/a1xnorb1 a1out_2 0.54fF
C1573 4bitadder_0/XOR_2/w_62_n20# 4bitadder_0/XOR_2/abar 0.02fF
C1574 comparator_0/t1 comparator_0/t2 0.18fF
C1575 gnd s0 8.09fF
C1576 enable_1/and_2/w_n43_8# a2 0.09fF
C1577 enable_1/and_4/w_26_9# b0out_1 0.03fF
C1578 s0 4bitadder_1/XOR_2/w_62_37# 0.13fF
C1579 enable_0/and_6/w_26_9# enable_0/and_6/a_n26_14# 0.09fF
C1580 4bitadder_1/fulladder_2/and_1/w_n43_8# a2out_1 0.09fF
C1581 enable_1/and_4/w_26_9# vdd 0.03fF
C1582 4bitadder_0/XOR_0/w_62_37# s0 0.13fF
C1583 4bitadder_0/XOR_0/abar 4bitadder_0/XOR_0/w_n34_n1# 0.03fF
C1584 4bitadder_0/XOR_1/out a1out_0 1.87fF
C1585 4bitadder_0/fulladder_1/and_1/w_26_9# 4bitadder_0/fulladder_1/or_0/b 0.03fF
C1586 enable_2/and_1/w_n43_8# enable_2/and_1/a_n26_14# 0.02fF
C1587 4bitadder_0/c2 4bitadder_0/fulladder_2/XOR_1/w_62_37# 0.13fF
C1588 out1 gnd 0.01fF
C1589 enable_1/and_5/w_n43_8# enable_1/en 0.09fF
C1590 vdd decoder_0/and_1/b 0.04fF
C1591 comparator_0/a1xnorb1 comparator_0/a0xnorb0 0.40fF
C1592 enable_2/en a0 0.27fF
C1593 4bitadder_0/fulladder_1/or_0/w_n48_101# 4bitadder_0/fulladder_1/or_0/a 0.12fF
C1594 4bitadder_0/fulladder_0/XOR_0/w_62_37# a0out_0 0.02fF
C1595 enable_2/en enable_2/and_3/w_n43_8# 0.09fF
C1596 4bitadder_1/XOR_0/w_16_n1# s0 0.11fF
C1597 b3out_2 b2out_2 0.43fF
C1598 comparator_0/5input_AND_1/not_0/in comparator_0/5input_AND_1/w_68_n82# 0.02fF
C1599 4bitadder_0/c2 s2_add 0.04fF
C1600 4bitadder_0/fulladder_1/XOR_1/w_n34_n1# vdd 0.02fF
C1601 enable_2/and_2/w_n43_8# vdd 0.07fF
C1602 4bitadder_1/fulladder_3/and_0/a_n26_14# 4bitadder_1/c3 0.10fF
C1603 4bitadder_0/fulladder_3/XOR_0/w_62_n20# 4bitadder_0/fulladder_3/XOR_0/abar 0.02fF
C1604 b1 enable_0/and_5/a_n26_14# 0.31fF
C1605 a0 a2 0.40fF
C1606 4bitadder_1/fulladder_3/axorb 4bitadder_1/fulladder_3/XOR_1/abar 0.13fF
C1607 4bitadder_0/fulladder_0/XOR_0/bbar 4bitadder_0/b0xorM 0.02fF
C1608 decoder_0/and_2/w_n43_8# decoder_0/and_2/a_n26_14# 0.02fF
C1609 4bitadder_1/fulladder_2/or_0/w_n48_101# 4bitadder_1/fulladder_2/or_0/a 0.12fF
C1610 comparator_0/5input_AND_1/w_106_n113# comparator_0/a3xnorb3 0.17fF
C1611 comparator_0/xnor_1/not_0/w_n2_10# comparator_0/xnor_1/not_0/in 0.09fF
C1612 vdd 4bitadder_1/fulladder_1/and_0/w_26_9# 0.03fF
C1613 vdd comparator_0/5input_AND_1/w_n37_15# 0.05fF
C1614 enable_1/and_7/a_n26_14# b3 0.31fF
C1615 vdd 4bitadder_1/c3 0.12fF
C1616 s0 decoder_0/not_0/w_n2_10# 0.09fF
C1617 gnd b1out_1 1.08fF
C1618 b3 a1 0.31fF
C1619 enable_3/en a2 0.25fF
C1620 4bitadder_1/fulladder_1/XOR_1/w_62_37# s1_sub 0.02fF
C1621 4bitadder_1/fulladder_1/axorb 4bitadder_1/fulladder_1/XOR_1/w_n34_n1# 0.11fF
C1622 4bitadder_0/fulladder_2/and_0/w_n43_8# vdd 0.07fF
C1623 comparator_0/b1bar comparator_0/4input_AND_1/not_0/in 0.18fF
C1624 a3out_2 comparator_0/and_0/w_n43_8# 0.09fF
C1625 vdd comparator_0/4input_OR_1/NOT_0/w_n2_10# 0.18fF
C1626 b2 b1 0.34fF
C1627 4bitadder_0/fulladder_0/XOR_1/w_16_n1# 4bitadder_0/fulladder_0/XOR_1/bbar 0.03fF
C1628 4bitadder_0/fulladder_0/XOR_1/w_62_n20# s0_add 0.04fF
C1629 4bitadder_0/fulladder_0/XOR_1/w_n34_n1# 4bitadder_0/fulladder_0/XOR_1/abar 0.03fF
C1630 4bitadder_0/XOR_1/abar b1out_0 0.13fF
C1631 enable_0/en vdd 0.93fF
C1632 a2out_2 b1out_2 1.07fF
C1633 b2out_2 a1out_2 0.65fF
C1634 4bitadder_0/XOR_1/w_62_37# s0 0.13fF
C1635 comparator_0/not_7/w_n2_10# comparator_0/a3bar 0.03fF
C1636 gnd b1out_0 0.52fF
C1637 comparator_0/xnor_3/XOR_0/w_62_n20# comparator_0/xnor_3/XOR_0/abar 0.02fF
C1638 4bitadder_0/fulladder_2/and_1/w_n43_8# a2out_0 0.09fF
C1639 comparator_0/3input_AND_1/not_0/in comparator_0/3input_AND_1/w_69_n71# 0.02fF
C1640 enable_0/en a3 0.37fF
C1641 4bitadder_0/fulladder_3/or_0/a vdd 0.14fF
C1642 4bitadder_0/fulladder_2/XOR_0/abar gnd 0.15fF
C1643 comparator_0/4input_OR_1/NOT_0/w_n2_10# bga 0.03fF
C1644 4bitadder_1/fulladder_0/XOR_1/w_62_n20# s0_sub 0.04fF
C1645 4bitadder_0/XOR_2/out s0 0.19fF
C1646 vdd equal 0.04fF
C1647 vdd enable_0/and_5/w_26_9# 0.03fF
C1648 decoder_0/and_3/a_n26_14# Gnd 0.05fF
C1649 s1 Gnd 1.48fF
C1650 decoder_0/and_3/w_26_9# Gnd 0.82fF
C1651 decoder_0/and_3/w_n43_8# Gnd 0.82fF
C1652 decoder_0/and_2/a_n26_14# Gnd 0.05fF
C1653 decoder_0/and_2/w_26_9# Gnd 0.82fF
C1654 decoder_0/and_2/w_n43_8# Gnd 0.82fF
C1655 decoder_0/and_1/a_n26_14# Gnd 0.05fF
C1656 decoder_0/and_1/w_26_9# Gnd 0.82fF
C1657 decoder_0/and_1/w_n43_8# Gnd 0.82fF
C1658 decoder_0/and_0/a_n26_14# Gnd 0.05fF
C1659 decoder_0/and_0/w_26_9# Gnd 0.82fF
C1660 decoder_0/and_0/w_n43_8# Gnd 0.82fF
C1661 decoder_0/not_1/w_n2_10# Gnd 0.90fF
C1662 decoder_0/not_0/w_n2_10# Gnd 0.90fF
C1663 4bitadder_1/XOR_3/abar Gnd 0.11fF
C1664 4bitadder_1/XOR_3/bbar Gnd 0.06fF
C1665 4bitadder_1/XOR_3/w_62_n20# Gnd 0.87fF
C1666 4bitadder_1/XOR_3/w_16_n1# Gnd 0.75fF
C1667 4bitadder_1/XOR_3/w_n34_n1# Gnd 0.75fF
C1668 4bitadder_1/XOR_3/w_62_37# Gnd 0.72fF
C1669 4bitadder_1/XOR_2/abar Gnd 0.11fF
C1670 4bitadder_1/XOR_2/bbar Gnd 0.06fF
C1671 4bitadder_1/XOR_2/w_62_n20# Gnd 0.87fF
C1672 4bitadder_1/XOR_2/w_16_n1# Gnd 0.75fF
C1673 4bitadder_1/XOR_2/w_n34_n1# Gnd 0.75fF
C1674 4bitadder_1/XOR_2/w_62_37# Gnd 0.72fF
C1675 4bitadder_1/XOR_1/abar Gnd 0.11fF
C1676 4bitadder_1/XOR_1/bbar Gnd 0.06fF
C1677 s0 Gnd 36.69fF
C1678 b1out_1 Gnd 3.47fF
C1679 4bitadder_1/XOR_1/w_62_n20# Gnd 0.87fF
C1680 4bitadder_1/XOR_1/w_16_n1# Gnd 0.75fF
C1681 4bitadder_1/XOR_1/w_n34_n1# Gnd 0.75fF
C1682 4bitadder_1/XOR_1/w_62_37# Gnd 0.72fF
C1683 4bitadder_1/XOR_0/abar Gnd 0.12fF
C1684 4bitadder_1/XOR_0/bbar Gnd 0.06fF
C1685 b0out_1 Gnd 3.02fF
C1686 4bitadder_1/XOR_0/w_62_n20# Gnd 0.87fF
C1687 4bitadder_1/XOR_0/w_16_n1# Gnd 0.75fF
C1688 4bitadder_1/XOR_0/w_n34_n1# Gnd 0.75fF
C1689 4bitadder_1/XOR_0/w_62_37# Gnd 0.72fF
C1690 4bitadder_1/fulladder_3/XOR_1/abar Gnd 0.11fF
C1691 4bitadder_1/fulladder_3/XOR_1/bbar Gnd 0.06fF
C1692 s3_sub Gnd 1.05fF
C1693 4bitadder_1/fulladder_3/XOR_1/w_62_n20# Gnd 0.87fF
C1694 4bitadder_1/fulladder_3/XOR_1/w_16_n1# Gnd 0.75fF
C1695 4bitadder_1/fulladder_3/XOR_1/w_n34_n1# Gnd 0.75fF
C1696 4bitadder_1/fulladder_3/XOR_1/w_62_37# Gnd 0.72fF
C1697 4bitadder_1/fulladder_3/or_0/b Gnd 2.26fF
C1698 4bitadder_1/fulladder_3/and_1/a_n26_14# Gnd 0.05fF
C1699 a3out_1 Gnd 7.67fF
C1700 4bitadder_1/fulladder_3/and_1/w_26_9# Gnd 0.82fF
C1701 4bitadder_1/fulladder_3/and_1/w_n43_8# Gnd 0.82fF
C1702 4bitadder_1/fulladder_3/XOR_0/abar Gnd 0.11fF
C1703 4bitadder_1/fulladder_3/XOR_0/bbar Gnd 0.06fF
C1704 4bitadder_1/fulladder_3/XOR_0/w_62_n20# Gnd 0.87fF
C1705 4bitadder_1/fulladder_3/XOR_0/w_16_n1# Gnd 0.75fF
C1706 4bitadder_1/fulladder_3/XOR_0/w_n34_n1# Gnd 0.75fF
C1707 4bitadder_1/fulladder_3/XOR_0/w_62_37# Gnd 0.72fF
C1708 4bitadder_1/fulladder_3/or_0/a Gnd 1.96fF
C1709 4bitadder_1/fulladder_3/and_0/a_n26_14# Gnd 0.05fF
C1710 4bitadder_1/c3 Gnd 2.24fF
C1711 4bitadder_1/fulladder_3/axorb Gnd 3.25fF
C1712 4bitadder_1/fulladder_3/and_0/w_26_9# Gnd 0.82fF
C1713 4bitadder_1/fulladder_3/and_0/w_n43_8# Gnd 0.82fF
C1714 fc_sub Gnd 0.60fF
C1715 4bitadder_1/fulladder_3/or_0/a_n15_32# Gnd 0.17fF
C1716 4bitadder_1/fulladder_3/or_0/w_58_101# Gnd 1.55fF
C1717 4bitadder_1/fulladder_3/or_0/w_n48_101# Gnd 2.56fF
C1718 4bitadder_1/fulladder_2/XOR_1/abar Gnd 0.11fF
C1719 4bitadder_1/fulladder_2/XOR_1/bbar Gnd 0.06fF
C1720 s2_sub Gnd 0.72fF
C1721 4bitadder_1/fulladder_2/XOR_1/w_62_n20# Gnd 0.87fF
C1722 4bitadder_1/fulladder_2/XOR_1/w_16_n1# Gnd 0.75fF
C1723 4bitadder_1/fulladder_2/XOR_1/w_n34_n1# Gnd 0.75fF
C1724 4bitadder_1/fulladder_2/XOR_1/w_62_37# Gnd 0.72fF
C1725 4bitadder_1/fulladder_2/or_0/b Gnd 2.26fF
C1726 4bitadder_1/fulladder_2/and_1/a_n26_14# Gnd 0.05fF
C1727 4bitadder_1/XOR_2/out Gnd 2.12fF
C1728 4bitadder_1/fulladder_2/and_1/w_26_9# Gnd 0.82fF
C1729 4bitadder_1/fulladder_2/and_1/w_n43_8# Gnd 0.82fF
C1730 4bitadder_1/fulladder_2/XOR_0/abar Gnd 0.11fF
C1731 4bitadder_1/fulladder_2/XOR_0/bbar Gnd 0.06fF
C1732 4bitadder_1/fulladder_2/XOR_0/w_62_n20# Gnd 0.87fF
C1733 4bitadder_1/fulladder_2/XOR_0/w_16_n1# Gnd 0.75fF
C1734 4bitadder_1/fulladder_2/XOR_0/w_n34_n1# Gnd 0.75fF
C1735 4bitadder_1/fulladder_2/XOR_0/w_62_37# Gnd 0.72fF
C1736 4bitadder_1/fulladder_2/or_0/a Gnd 1.96fF
C1737 4bitadder_1/fulladder_2/and_0/a_n26_14# Gnd 0.05fF
C1738 4bitadder_1/fulladder_2/axorb Gnd 3.25fF
C1739 4bitadder_1/fulladder_2/and_0/w_26_9# Gnd 0.82fF
C1740 4bitadder_1/fulladder_2/and_0/w_n43_8# Gnd 0.82fF
C1741 4bitadder_1/fulladder_2/or_0/a_n15_32# Gnd 0.17fF
C1742 4bitadder_1/fulladder_2/or_0/w_58_101# Gnd 1.55fF
C1743 4bitadder_1/fulladder_2/or_0/w_n48_101# Gnd 2.56fF
C1744 4bitadder_1/fulladder_1/XOR_1/abar Gnd 0.11fF
C1745 4bitadder_1/fulladder_1/XOR_1/bbar Gnd 0.06fF
C1746 s1_sub Gnd 1.01fF
C1747 4bitadder_1/fulladder_1/XOR_1/w_62_n20# Gnd 0.87fF
C1748 4bitadder_1/fulladder_1/XOR_1/w_16_n1# Gnd 0.75fF
C1749 4bitadder_1/fulladder_1/XOR_1/w_n34_n1# Gnd 0.75fF
C1750 4bitadder_1/fulladder_1/XOR_1/w_62_37# Gnd 0.72fF
C1751 4bitadder_1/fulladder_1/or_0/b Gnd 2.26fF
C1752 4bitadder_1/fulladder_1/and_1/a_n26_14# Gnd 0.05fF
C1753 4bitadder_1/XOR_1/out Gnd 2.08fF
C1754 4bitadder_1/fulladder_1/and_1/w_26_9# Gnd 0.82fF
C1755 4bitadder_1/fulladder_1/and_1/w_n43_8# Gnd 0.82fF
C1756 4bitadder_1/fulladder_1/XOR_0/abar Gnd 0.11fF
C1757 4bitadder_1/fulladder_1/XOR_0/bbar Gnd 0.06fF
C1758 4bitadder_1/fulladder_1/XOR_0/w_62_n20# Gnd 0.87fF
C1759 4bitadder_1/fulladder_1/XOR_0/w_16_n1# Gnd 0.75fF
C1760 4bitadder_1/fulladder_1/XOR_0/w_n34_n1# Gnd 0.75fF
C1761 4bitadder_1/fulladder_1/XOR_0/w_62_37# Gnd 0.72fF
C1762 4bitadder_1/fulladder_1/or_0/a Gnd 1.96fF
C1763 4bitadder_1/fulladder_1/and_0/a_n26_14# Gnd 0.05fF
C1764 4bitadder_1/fulladder_1/axorb Gnd 3.25fF
C1765 4bitadder_1/fulladder_1/and_0/w_26_9# Gnd 0.82fF
C1766 4bitadder_1/fulladder_1/and_0/w_n43_8# Gnd 0.82fF
C1767 4bitadder_1/fulladder_1/or_0/a_n15_32# Gnd 0.17fF
C1768 4bitadder_1/fulladder_1/or_0/w_58_101# Gnd 1.55fF
C1769 4bitadder_1/fulladder_1/or_0/w_n48_101# Gnd 2.56fF
C1770 4bitadder_1/fulladder_0/XOR_1/abar Gnd 0.11fF
C1771 4bitadder_1/fulladder_0/XOR_1/bbar Gnd 0.06fF
C1772 s0_sub Gnd 0.46fF
C1773 4bitadder_1/fulladder_0/XOR_1/w_62_n20# Gnd 0.87fF
C1774 4bitadder_1/fulladder_0/XOR_1/w_16_n1# Gnd 0.75fF
C1775 4bitadder_1/fulladder_0/XOR_1/w_n34_n1# Gnd 0.75fF
C1776 4bitadder_1/fulladder_0/XOR_1/w_62_37# Gnd 0.72fF
C1777 4bitadder_1/fulladder_0/or_0/b Gnd 2.26fF
C1778 4bitadder_1/fulladder_0/and_1/a_n26_14# Gnd 0.05fF
C1779 a0_out1 Gnd 7.61fF
C1780 4bitadder_1/b0xorM Gnd 2.11fF
C1781 4bitadder_1/fulladder_0/and_1/w_26_9# Gnd 0.82fF
C1782 4bitadder_1/fulladder_0/and_1/w_n43_8# Gnd 0.82fF
C1783 4bitadder_1/fulladder_0/XOR_0/abar Gnd 0.11fF
C1784 4bitadder_1/fulladder_0/XOR_0/bbar Gnd 0.06fF
C1785 4bitadder_1/fulladder_0/XOR_0/w_62_n20# Gnd 0.87fF
C1786 4bitadder_1/fulladder_0/XOR_0/w_16_n1# Gnd 0.75fF
C1787 4bitadder_1/fulladder_0/XOR_0/w_n34_n1# Gnd 0.75fF
C1788 4bitadder_1/fulladder_0/XOR_0/w_62_37# Gnd 0.72fF
C1789 4bitadder_1/fulladder_0/or_0/a Gnd 1.96fF
C1790 4bitadder_1/fulladder_0/and_0/a_n26_14# Gnd 0.05fF
C1791 4bitadder_1/fulladder_0/axorb Gnd 3.25fF
C1792 4bitadder_1/fulladder_0/and_0/w_26_9# Gnd 0.82fF
C1793 4bitadder_1/fulladder_0/and_0/w_n43_8# Gnd 0.82fF
C1794 4bitadder_1/fulladder_0/or_0/a_n15_32# Gnd 0.17fF
C1795 4bitadder_1/fulladder_0/or_0/w_58_101# Gnd 1.55fF
C1796 4bitadder_1/fulladder_0/or_0/w_n48_101# Gnd 2.56fF
C1797 comparator_0/a2bar Gnd 5.34fF
C1798 comparator_0/3input_AND_1/w_69_n71# Gnd 1.13fF
C1799 comparator_0/3input_AND_1/w_32_n21# Gnd 1.13fF
C1800 comparator_0/3input_AND_1/w_n14_24# Gnd 1.13fF
C1801 gnd Gnd 99.11fF
C1802 comparator_0/t2 Gnd 3.00fF
C1803 comparator_0/3input_AND_1/not_0/in Gnd 1.59fF
C1804 comparator_0/3input_AND_1/not_0/w_n2_10# Gnd 0.90fF
C1805 comparator_0/b2bar Gnd 5.92fF
C1806 comparator_0/3input_AND_0/w_69_n71# Gnd 1.13fF
C1807 comparator_0/3input_AND_0/w_32_n21# Gnd 1.13fF
C1808 comparator_0/3input_AND_0/w_n14_24# Gnd 1.13fF
C1809 comparator_0/t6 Gnd 2.94fF
C1810 comparator_0/3input_AND_0/not_0/in Gnd 1.59fF
C1811 comparator_0/3input_AND_0/not_0/w_n2_10# Gnd 0.90fF
C1812 comparator_0/a2xnorb2 Gnd 18.99fF
C1813 comparator_0/4input_AND_2/w_68_n95# Gnd 1.13fF
C1814 comparator_0/4input_AND_2/w_29_n46# Gnd 1.13fF
C1815 comparator_0/4input_AND_2/w_n8_2# Gnd 1.13fF
C1816 comparator_0/4input_AND_2/w_n47_52# Gnd 1.13fF
C1817 comparator_0/t3 Gnd 4.44fF
C1818 comparator_0/4input_AND_2/not_0/in Gnd 2.38fF
C1819 comparator_0/4input_AND_2/not_0/w_n2_10# Gnd 0.90fF
C1820 comparator_0/and_1/a_n26_14# Gnd 0.05fF
C1821 comparator_0/a3bar Gnd 4.39fF
C1822 comparator_0/and_1/w_26_9# Gnd 0.82fF
C1823 comparator_0/and_1/w_n43_8# Gnd 0.82fF
C1824 comparator_0/4input_AND_1/w_68_n95# Gnd 1.13fF
C1825 comparator_0/4input_AND_1/w_29_n46# Gnd 1.13fF
C1826 comparator_0/4input_AND_1/w_n8_2# Gnd 1.13fF
C1827 comparator_0/4input_AND_1/w_n47_52# Gnd 1.13fF
C1828 comparator_0/t7 Gnd 4.39fF
C1829 comparator_0/4input_AND_1/not_0/in Gnd 2.38fF
C1830 comparator_0/4input_AND_1/not_0/w_n2_10# Gnd 0.90fF
C1831 comparator_0/4input_AND_0/w_68_n95# Gnd 1.13fF
C1832 comparator_0/4input_AND_0/w_29_n46# Gnd 1.13fF
C1833 comparator_0/4input_AND_0/w_n8_2# Gnd 1.13fF
C1834 comparator_0/4input_AND_0/w_n47_52# Gnd 1.13fF
C1835 equal Gnd 0.23fF
C1836 comparator_0/4input_AND_0/not_0/in Gnd 2.38fF
C1837 comparator_0/4input_AND_0/not_0/w_n2_10# Gnd 0.90fF
C1838 comparator_0/and_0/a_n26_14# Gnd 0.05fF
C1839 comparator_0/b3bar Gnd 0.68fF
C1840 comparator_0/and_0/w_26_9# Gnd 0.82fF
C1841 comparator_0/and_0/w_n43_8# Gnd 0.82fF
C1842 comparator_0/5input_AND_1/w_106_n113# Gnd 0.81fF
C1843 comparator_0/5input_AND_1/w_68_n82# Gnd 0.81fF
C1844 comparator_0/5input_AND_1/w_31_n55# Gnd 1.18fF
C1845 comparator_0/5input_AND_1/w_n4_n20# Gnd 0.89fF
C1846 comparator_0/5input_AND_1/w_n37_15# Gnd 0.89fF
C1847 comparator_0/t4 Gnd 2.77fF
C1848 comparator_0/5input_AND_1/not_0/in Gnd 2.73fF
C1849 comparator_0/5input_AND_1/not_0/w_n2_10# Gnd 0.90fF
C1850 comparator_0/5input_AND_0/w_106_n113# Gnd 0.81fF
C1851 comparator_0/5input_AND_0/w_68_n82# Gnd 0.81fF
C1852 comparator_0/5input_AND_0/w_31_n55# Gnd 1.18fF
C1853 comparator_0/5input_AND_0/w_n4_n20# Gnd 0.89fF
C1854 comparator_0/5input_AND_0/w_n37_15# Gnd 0.89fF
C1855 comparator_0/t8 Gnd 1.96fF
C1856 comparator_0/5input_AND_0/not_0/in Gnd 2.73fF
C1857 comparator_0/5input_AND_0/not_0/w_n2_10# Gnd 0.90fF
C1858 comparator_0/not_7/w_n2_10# Gnd 0.90fF
C1859 comparator_0/not_6/w_n2_10# Gnd 0.90fF
C1860 comparator_0/a1bar Gnd 5.03fF
C1861 comparator_0/not_5/w_n2_10# Gnd 0.90fF
C1862 comparator_0/xnor_3/XOR_0/abar Gnd 0.11fF
C1863 comparator_0/xnor_3/XOR_0/bbar Gnd 0.06fF
C1864 comparator_0/xnor_3/not_0/in Gnd 0.39fF
C1865 boout_2 Gnd 8.80fF
C1866 a0out_2 Gnd 32.03fF
C1867 comparator_0/xnor_3/XOR_0/w_62_n20# Gnd 0.87fF
C1868 comparator_0/xnor_3/XOR_0/w_16_n1# Gnd 0.75fF
C1869 comparator_0/xnor_3/XOR_0/w_n34_n1# Gnd 0.75fF
C1870 comparator_0/xnor_3/XOR_0/w_62_37# Gnd 0.72fF
C1871 comparator_0/a0xnorb0 Gnd 2.96fF
C1872 comparator_0/xnor_3/not_0/w_n2_10# Gnd 0.90fF
C1873 comparator_0/xnor_2/XOR_0/abar Gnd 0.11fF
C1874 comparator_0/xnor_2/XOR_0/bbar Gnd 0.06fF
C1875 comparator_0/xnor_2/not_0/in Gnd 0.39fF
C1876 b1out_2 Gnd 55.09fF
C1877 a1out_2 Gnd 41.81fF
C1878 comparator_0/xnor_2/XOR_0/w_62_n20# Gnd 0.87fF
C1879 comparator_0/xnor_2/XOR_0/w_16_n1# Gnd 0.75fF
C1880 comparator_0/xnor_2/XOR_0/w_n34_n1# Gnd 0.75fF
C1881 comparator_0/xnor_2/XOR_0/w_62_37# Gnd 0.72fF
C1882 comparator_0/xnor_2/not_0/w_n2_10# Gnd 0.90fF
C1883 comparator_0/4input_OR_1/w_n58_n43# Gnd 2.55fF
C1884 bga Gnd 0.14fF
C1885 comparator_0/4input_OR_1/y Gnd 1.46fF
C1886 comparator_0/4input_OR_1/NOT_0/w_n2_10# Gnd 0.90fF
C1887 comparator_0/a0bar Gnd 6.16fF
C1888 comparator_0/not_4/w_n2_10# Gnd 0.90fF
C1889 comparator_0/xnor_1/XOR_0/abar Gnd 0.11fF
C1890 comparator_0/xnor_1/XOR_0/bbar Gnd 0.06fF
C1891 comparator_0/xnor_1/not_0/in Gnd 0.39fF
C1892 b2out_2 Gnd 46.65fF
C1893 a2out_2 Gnd 27.86fF
C1894 comparator_0/xnor_1/XOR_0/w_62_n20# Gnd 0.87fF
C1895 comparator_0/xnor_1/XOR_0/w_16_n1# Gnd 0.75fF
C1896 comparator_0/xnor_1/XOR_0/w_n34_n1# Gnd 0.75fF
C1897 comparator_0/xnor_1/XOR_0/w_62_37# Gnd 0.72fF
C1898 comparator_0/xnor_1/not_0/w_n2_10# Gnd 0.90fF
C1899 comparator_0/not_3/w_n2_10# Gnd 0.90fF
C1900 comparator_0/xnor_0/XOR_0/abar Gnd 0.11fF
C1901 comparator_0/xnor_0/XOR_0/bbar Gnd 0.06fF
C1902 comparator_0/xnor_0/not_0/in Gnd 0.39fF
C1903 b3out_2 Gnd 29.74fF
C1904 a3out_2 Gnd 20.89fF
C1905 comparator_0/xnor_0/XOR_0/w_62_n20# Gnd 0.87fF
C1906 comparator_0/xnor_0/XOR_0/w_16_n1# Gnd 0.75fF
C1907 comparator_0/xnor_0/XOR_0/w_n34_n1# Gnd 0.75fF
C1908 comparator_0/xnor_0/XOR_0/w_62_37# Gnd 0.72fF
C1909 comparator_0/xnor_0/not_0/w_n2_10# Gnd 0.90fF
C1910 comparator_0/not_2/w_n2_10# Gnd 0.90fF
C1911 comparator_0/4input_OR_0/w_n58_n43# Gnd 2.55fF
C1912 agb Gnd 0.14fF
C1913 comparator_0/4input_OR_0/y Gnd 1.46fF
C1914 vdd Gnd 121.02fF
C1915 comparator_0/4input_OR_0/NOT_0/w_n2_10# Gnd 0.90fF
C1916 comparator_0/b1bar Gnd 4.66fF
C1917 comparator_0/not_1/w_n2_10# Gnd 0.90fF
C1918 comparator_0/b0bar Gnd 6.97fF
C1919 comparator_0/not_0/w_n2_10# Gnd 0.90fF
C1920 4bitadder_0/XOR_3/abar Gnd 0.11fF
C1921 4bitadder_0/XOR_3/bbar Gnd 0.06fF
C1922 4bitadder_0/XOR_3/w_62_n20# Gnd 0.87fF
C1923 4bitadder_0/XOR_3/w_16_n1# Gnd 0.75fF
C1924 4bitadder_0/XOR_3/w_n34_n1# Gnd 0.75fF
C1925 4bitadder_0/XOR_3/w_62_37# Gnd 0.72fF
C1926 4bitadder_0/XOR_2/abar Gnd 0.11fF
C1927 4bitadder_0/XOR_2/bbar Gnd 0.06fF
C1928 4bitadder_0/XOR_2/w_62_n20# Gnd 0.87fF
C1929 4bitadder_0/XOR_2/w_16_n1# Gnd 0.75fF
C1930 4bitadder_0/XOR_2/w_n34_n1# Gnd 0.75fF
C1931 4bitadder_0/XOR_2/w_62_37# Gnd 0.72fF
C1932 4bitadder_0/XOR_1/abar Gnd 0.11fF
C1933 4bitadder_0/XOR_1/bbar Gnd 0.06fF
C1934 4bitadder_0/XOR_1/w_62_n20# Gnd 0.87fF
C1935 4bitadder_0/XOR_1/w_16_n1# Gnd 0.75fF
C1936 4bitadder_0/XOR_1/w_n34_n1# Gnd 0.75fF
C1937 4bitadder_0/XOR_1/w_62_37# Gnd 0.72fF
C1938 4bitadder_0/XOR_0/abar Gnd 0.12fF
C1939 4bitadder_0/XOR_0/bbar Gnd 0.06fF
C1940 4bitadder_0/XOR_0/w_62_n20# Gnd 0.87fF
C1941 4bitadder_0/XOR_0/w_16_n1# Gnd 0.75fF
C1942 4bitadder_0/XOR_0/w_n34_n1# Gnd 0.75fF
C1943 4bitadder_0/XOR_0/w_62_37# Gnd 0.72fF
C1944 4bitadder_0/fulladder_3/XOR_1/abar Gnd 0.11fF
C1945 4bitadder_0/fulladder_3/XOR_1/bbar Gnd 0.06fF
C1946 s3_add Gnd 0.74fF
C1947 4bitadder_0/fulladder_3/XOR_1/w_62_n20# Gnd 0.87fF
C1948 4bitadder_0/fulladder_3/XOR_1/w_16_n1# Gnd 0.75fF
C1949 4bitadder_0/fulladder_3/XOR_1/w_n34_n1# Gnd 0.75fF
C1950 4bitadder_0/fulladder_3/XOR_1/w_62_37# Gnd 0.72fF
C1951 4bitadder_0/fulladder_3/or_0/b Gnd 2.26fF
C1952 4bitadder_0/fulladder_3/and_1/a_n26_14# Gnd 0.05fF
C1953 a3out_0 Gnd 7.66fF
C1954 4bitadder_0/fulladder_3/and_1/w_26_9# Gnd 0.82fF
C1955 4bitadder_0/fulladder_3/and_1/w_n43_8# Gnd 0.82fF
C1956 4bitadder_0/fulladder_3/XOR_0/abar Gnd 0.11fF
C1957 4bitadder_0/fulladder_3/XOR_0/bbar Gnd 0.06fF
C1958 4bitadder_0/fulladder_3/XOR_0/w_62_n20# Gnd 0.87fF
C1959 4bitadder_0/fulladder_3/XOR_0/w_16_n1# Gnd 0.75fF
C1960 4bitadder_0/fulladder_3/XOR_0/w_n34_n1# Gnd 0.75fF
C1961 4bitadder_0/fulladder_3/XOR_0/w_62_37# Gnd 0.72fF
C1962 4bitadder_0/fulladder_3/or_0/a Gnd 1.96fF
C1963 4bitadder_0/fulladder_3/and_0/a_n26_14# Gnd 0.05fF
C1964 4bitadder_0/c3 Gnd 2.24fF
C1965 4bitadder_0/fulladder_3/axorb Gnd 3.25fF
C1966 4bitadder_0/fulladder_3/and_0/w_26_9# Gnd 0.82fF
C1967 4bitadder_0/fulladder_3/and_0/w_n43_8# Gnd 0.82fF
C1968 fc_add Gnd 0.54fF
C1969 4bitadder_0/fulladder_3/or_0/a_n15_32# Gnd 0.17fF
C1970 4bitadder_0/fulladder_3/or_0/w_58_101# Gnd 1.55fF
C1971 4bitadder_0/fulladder_3/or_0/w_n48_101# Gnd 2.56fF
C1972 4bitadder_0/fulladder_2/XOR_1/abar Gnd 0.11fF
C1973 4bitadder_0/fulladder_2/XOR_1/bbar Gnd 0.06fF
C1974 s2_add Gnd 0.65fF
C1975 4bitadder_0/fulladder_2/XOR_1/w_62_n20# Gnd 0.87fF
C1976 4bitadder_0/fulladder_2/XOR_1/w_16_n1# Gnd 0.75fF
C1977 4bitadder_0/fulladder_2/XOR_1/w_n34_n1# Gnd 0.75fF
C1978 4bitadder_0/fulladder_2/XOR_1/w_62_37# Gnd 0.72fF
C1979 4bitadder_0/fulladder_2/or_0/b Gnd 2.26fF
C1980 4bitadder_0/fulladder_2/and_1/a_n26_14# Gnd 0.05fF
C1981 a2out_0 Gnd 7.81fF
C1982 4bitadder_0/XOR_2/out Gnd 2.12fF
C1983 4bitadder_0/fulladder_2/and_1/w_26_9# Gnd 0.82fF
C1984 4bitadder_0/fulladder_2/and_1/w_n43_8# Gnd 0.82fF
C1985 4bitadder_0/fulladder_2/XOR_0/abar Gnd 0.11fF
C1986 4bitadder_0/fulladder_2/XOR_0/bbar Gnd 0.06fF
C1987 4bitadder_0/fulladder_2/XOR_0/w_62_n20# Gnd 0.87fF
C1988 4bitadder_0/fulladder_2/XOR_0/w_16_n1# Gnd 0.75fF
C1989 4bitadder_0/fulladder_2/XOR_0/w_n34_n1# Gnd 0.75fF
C1990 4bitadder_0/fulladder_2/XOR_0/w_62_37# Gnd 0.72fF
C1991 4bitadder_0/fulladder_2/or_0/a Gnd 1.96fF
C1992 4bitadder_0/fulladder_2/and_0/a_n26_14# Gnd 0.05fF
C1993 4bitadder_0/fulladder_2/axorb Gnd 3.25fF
C1994 4bitadder_0/fulladder_2/and_0/w_26_9# Gnd 0.82fF
C1995 4bitadder_0/fulladder_2/and_0/w_n43_8# Gnd 0.82fF
C1996 4bitadder_0/fulladder_2/or_0/a_n15_32# Gnd 0.17fF
C1997 4bitadder_0/fulladder_2/or_0/w_58_101# Gnd 1.55fF
C1998 4bitadder_0/fulladder_2/or_0/w_n48_101# Gnd 2.56fF
C1999 4bitadder_0/fulladder_1/XOR_1/abar Gnd 0.11fF
C2000 4bitadder_0/fulladder_1/XOR_1/bbar Gnd 0.06fF
C2001 s1_add Gnd 1.15fF
C2002 4bitadder_0/fulladder_1/XOR_1/w_62_n20# Gnd 0.87fF
C2003 4bitadder_0/fulladder_1/XOR_1/w_16_n1# Gnd 0.75fF
C2004 4bitadder_0/fulladder_1/XOR_1/w_n34_n1# Gnd 0.75fF
C2005 4bitadder_0/fulladder_1/XOR_1/w_62_37# Gnd 0.72fF
C2006 4bitadder_0/fulladder_1/or_0/b Gnd 2.26fF
C2007 4bitadder_0/fulladder_1/and_1/a_n26_14# Gnd 0.05fF
C2008 a1out_0 Gnd 7.72fF
C2009 4bitadder_0/XOR_1/out Gnd 2.08fF
C2010 4bitadder_0/fulladder_1/and_1/w_26_9# Gnd 0.82fF
C2011 4bitadder_0/fulladder_1/and_1/w_n43_8# Gnd 0.82fF
C2012 4bitadder_0/fulladder_1/XOR_0/abar Gnd 0.11fF
C2013 4bitadder_0/fulladder_1/XOR_0/bbar Gnd 0.06fF
C2014 4bitadder_0/fulladder_1/XOR_0/w_62_n20# Gnd 0.87fF
C2015 4bitadder_0/fulladder_1/XOR_0/w_16_n1# Gnd 0.75fF
C2016 4bitadder_0/fulladder_1/XOR_0/w_n34_n1# Gnd 0.75fF
C2017 4bitadder_0/fulladder_1/XOR_0/w_62_37# Gnd 0.72fF
C2018 4bitadder_0/fulladder_1/or_0/a Gnd 1.96fF
C2019 4bitadder_0/fulladder_1/and_0/a_n26_14# Gnd 0.05fF
C2020 4bitadder_0/fulladder_1/axorb Gnd 3.25fF
C2021 4bitadder_0/fulladder_1/and_0/w_26_9# Gnd 0.82fF
C2022 4bitadder_0/fulladder_1/and_0/w_n43_8# Gnd 0.82fF
C2023 4bitadder_0/fulladder_1/or_0/a_n15_32# Gnd 0.17fF
C2024 4bitadder_0/fulladder_1/or_0/w_58_101# Gnd 1.55fF
C2025 4bitadder_0/fulladder_1/or_0/w_n48_101# Gnd 2.56fF
C2026 4bitadder_0/fulladder_0/XOR_1/abar Gnd 0.11fF
C2027 4bitadder_0/fulladder_0/XOR_1/bbar Gnd 0.06fF
C2028 s0_add Gnd 0.87fF
C2029 4bitadder_0/fulladder_0/XOR_1/w_62_n20# Gnd 0.87fF
C2030 4bitadder_0/fulladder_0/XOR_1/w_16_n1# Gnd 0.75fF
C2031 4bitadder_0/fulladder_0/XOR_1/w_n34_n1# Gnd 0.75fF
C2032 4bitadder_0/fulladder_0/XOR_1/w_62_37# Gnd 0.72fF
C2033 4bitadder_0/fulladder_0/or_0/b Gnd 2.26fF
C2034 4bitadder_0/fulladder_0/and_1/a_n26_14# Gnd 0.05fF
C2035 a0out_0 Gnd 7.55fF
C2036 4bitadder_0/b0xorM Gnd 2.11fF
C2037 4bitadder_0/fulladder_0/and_1/w_26_9# Gnd 0.82fF
C2038 4bitadder_0/fulladder_0/and_1/w_n43_8# Gnd 0.82fF
C2039 4bitadder_0/fulladder_0/XOR_0/abar Gnd 0.11fF
C2040 4bitadder_0/fulladder_0/XOR_0/bbar Gnd 0.06fF
C2041 4bitadder_0/fulladder_0/XOR_0/w_62_n20# Gnd 0.87fF
C2042 4bitadder_0/fulladder_0/XOR_0/w_16_n1# Gnd 0.75fF
C2043 4bitadder_0/fulladder_0/XOR_0/w_n34_n1# Gnd 0.75fF
C2044 4bitadder_0/fulladder_0/XOR_0/w_62_37# Gnd 0.72fF
C2045 4bitadder_0/fulladder_0/or_0/a Gnd 1.96fF
C2046 4bitadder_0/fulladder_0/and_0/a_n26_14# Gnd 0.05fF
C2047 4bitadder_0/fulladder_0/axorb Gnd 3.25fF
C2048 4bitadder_0/fulladder_0/and_0/w_26_9# Gnd 0.82fF
C2049 4bitadder_0/fulladder_0/and_0/w_n43_8# Gnd 0.82fF
C2050 4bitadder_0/fulladder_0/or_0/a_n15_32# Gnd 0.17fF
C2051 4bitadder_0/fulladder_0/or_0/w_58_101# Gnd 1.55fF
C2052 4bitadder_0/fulladder_0/or_0/w_n48_101# Gnd 2.56fF
C2053 out3 Gnd 0.20fF
C2054 AND_Block_0/and_3/a_n26_14# Gnd 0.05fF
C2055 b3out_3 Gnd 0.73fF
C2056 a3out_3 Gnd 0.75fF
C2057 AND_Block_0/and_3/w_26_9# Gnd 0.82fF
C2058 AND_Block_0/and_3/w_n43_8# Gnd 0.82fF
C2059 out2 Gnd 0.20fF
C2060 AND_Block_0/and_2/a_n26_14# Gnd 0.05fF
C2061 b2out_3 Gnd 0.74fF
C2062 a2out_3 Gnd 0.77fF
C2063 AND_Block_0/and_2/w_26_9# Gnd 0.82fF
C2064 AND_Block_0/and_2/w_n43_8# Gnd 0.82fF
C2065 out1 Gnd 0.21fF
C2066 AND_Block_0/and_1/a_n26_14# Gnd 0.05fF
C2067 b1out_3 Gnd 0.75fF
C2068 a1out_3 Gnd 0.79fF
C2069 AND_Block_0/and_1/w_26_9# Gnd 0.82fF
C2070 AND_Block_0/and_1/w_n43_8# Gnd 0.82fF
C2071 out0 Gnd 0.20fF
C2072 AND_Block_0/and_0/a_n26_14# Gnd 0.05fF
C2073 b0out_3 Gnd 0.72fF
C2074 AND_Block_0/and_0/w_26_9# Gnd 0.82fF
C2075 AND_Block_0/and_0/w_n43_8# Gnd 0.82fF
C2076 enable_3/and_4/a_n26_14# Gnd 0.05fF
C2077 b0 Gnd 1.59fF
C2078 enable_3/and_4/w_26_9# Gnd 0.82fF
C2079 enable_3/and_4/w_n43_8# Gnd 0.82fF
C2080 enable_3/and_3/a_n26_14# Gnd 0.05fF
C2081 a3 Gnd 1.58fF
C2082 enable_3/and_3/w_26_9# Gnd 0.82fF
C2083 enable_3/and_3/w_n43_8# Gnd 0.82fF
C2084 enable_3/and_2/a_n26_14# Gnd 0.05fF
C2085 a2 Gnd 1.49fF
C2086 enable_3/and_2/w_26_9# Gnd 0.82fF
C2087 enable_3/and_2/w_n43_8# Gnd 0.82fF
C2088 enable_3/and_1/a_n26_14# Gnd 0.05fF
C2089 enable_3/and_1/w_26_9# Gnd 0.82fF
C2090 enable_3/and_1/w_n43_8# Gnd 0.82fF
C2091 enable_3/and_0/a_n26_14# Gnd 0.05fF
C2092 a0 Gnd 1.49fF
C2093 enable_3/and_0/w_26_9# Gnd 0.82fF
C2094 enable_3/and_0/w_n43_8# Gnd 0.82fF
C2095 enable_3/and_6/a_n26_14# Gnd 0.05fF
C2096 b2 Gnd 1.57fF
C2097 enable_3/and_6/w_26_9# Gnd 0.82fF
C2098 enable_3/and_6/w_n43_8# Gnd 0.82fF
C2099 enable_3/and_7/a_n26_14# Gnd 0.05fF
C2100 b3 Gnd 1.60fF
C2101 enable_3/en Gnd 7.29fF
C2102 enable_3/and_7/w_26_9# Gnd 0.82fF
C2103 enable_3/and_7/w_n43_8# Gnd 0.82fF
C2104 enable_3/and_5/a_n26_14# Gnd 0.05fF
C2105 b1 Gnd 1.48fF
C2106 enable_3/and_5/w_26_9# Gnd 0.82fF
C2107 enable_3/and_5/w_n43_8# Gnd 0.82fF
C2108 enable_2/and_4/a_n26_14# Gnd 0.05fF
C2109 enable_2/and_4/w_26_9# Gnd 0.82fF
C2110 enable_2/and_4/w_n43_8# Gnd 0.82fF
C2111 enable_2/and_3/a_n26_14# Gnd 0.05fF
C2112 enable_2/and_3/w_26_9# Gnd 0.82fF
C2113 enable_2/and_3/w_n43_8# Gnd 0.82fF
C2114 enable_2/and_2/a_n26_14# Gnd 0.05fF
C2115 enable_2/and_2/w_26_9# Gnd 0.82fF
C2116 enable_2/and_2/w_n43_8# Gnd 0.82fF
C2117 enable_2/and_1/a_n26_14# Gnd 0.05fF
C2118 enable_2/and_1/w_26_9# Gnd 0.82fF
C2119 enable_2/and_1/w_n43_8# Gnd 0.82fF
C2120 enable_2/and_0/a_n26_14# Gnd 0.05fF
C2121 enable_2/and_0/w_26_9# Gnd 0.82fF
C2122 enable_2/and_0/w_n43_8# Gnd 0.82fF
C2123 enable_2/and_6/a_n26_14# Gnd 0.05fF
C2124 enable_2/and_6/w_26_9# Gnd 0.82fF
C2125 enable_2/and_6/w_n43_8# Gnd 0.82fF
C2126 enable_2/and_7/a_n26_14# Gnd 0.05fF
C2127 enable_2/en Gnd 2.76fF
C2128 enable_2/and_7/w_26_9# Gnd 0.82fF
C2129 enable_2/and_7/w_n43_8# Gnd 0.82fF
C2130 enable_2/and_5/a_n26_14# Gnd 0.05fF
C2131 enable_2/and_5/w_26_9# Gnd 0.82fF
C2132 enable_2/and_5/w_n43_8# Gnd 0.82fF
C2133 enable_1/and_4/a_n26_14# Gnd 0.05fF
C2134 enable_1/and_4/w_26_9# Gnd 0.82fF
C2135 enable_1/and_4/w_n43_8# Gnd 0.82fF
C2136 enable_1/and_3/a_n26_14# Gnd 0.05fF
C2137 enable_1/and_3/w_26_9# Gnd 0.82fF
C2138 enable_1/and_3/w_n43_8# Gnd 0.82fF
C2139 enable_1/and_2/a_n26_14# Gnd 0.05fF
C2140 enable_1/and_2/w_26_9# Gnd 0.82fF
C2141 enable_1/and_2/w_n43_8# Gnd 0.82fF
C2142 enable_1/and_1/a_n26_14# Gnd 0.05fF
C2143 enable_1/and_1/w_26_9# Gnd 0.82fF
C2144 enable_1/and_1/w_n43_8# Gnd 0.82fF
C2145 enable_1/and_0/a_n26_14# Gnd 0.05fF
C2146 enable_1/and_0/w_26_9# Gnd 0.82fF
C2147 enable_1/and_0/w_n43_8# Gnd 0.82fF
C2148 enable_1/and_6/a_n26_14# Gnd 0.05fF
C2149 enable_1/and_6/w_26_9# Gnd 0.82fF
C2150 enable_1/and_6/w_n43_8# Gnd 0.82fF
C2151 enable_1/and_7/a_n26_14# Gnd 0.05fF
C2152 enable_1/en Gnd 2.89fF
C2153 enable_1/and_7/w_26_9# Gnd 0.82fF
C2154 enable_1/and_7/w_n43_8# Gnd 0.82fF
C2155 enable_1/and_5/a_n26_14# Gnd 0.05fF
C2156 enable_1/and_5/w_26_9# Gnd 0.82fF
C2157 enable_1/and_5/w_n43_8# Gnd 0.82fF
C2158 b0out_0 Gnd 3.00fF
C2159 enable_0/and_4/a_n26_14# Gnd 0.05fF
C2160 enable_0/and_4/w_26_9# Gnd 0.82fF
C2161 enable_0/and_4/w_n43_8# Gnd 0.82fF
C2162 enable_0/and_3/a_n26_14# Gnd 0.05fF
C2163 enable_0/and_3/w_26_9# Gnd 0.82fF
C2164 enable_0/and_3/w_n43_8# Gnd 0.82fF
C2165 enable_0/and_2/a_n26_14# Gnd 0.05fF
C2166 enable_0/and_2/w_26_9# Gnd 0.82fF
C2167 enable_0/and_2/w_n43_8# Gnd 0.82fF
C2168 enable_0/and_1/a_n26_14# Gnd 0.05fF
C2169 enable_0/and_1/w_26_9# Gnd 0.82fF
C2170 enable_0/and_1/w_n43_8# Gnd 0.82fF
C2171 enable_0/and_0/a_n26_14# Gnd 0.05fF
C2172 enable_0/and_0/w_26_9# Gnd 0.82fF
C2173 enable_0/and_0/w_n43_8# Gnd 0.82fF
C2174 enable_0/and_6/a_n26_14# Gnd 0.05fF
C2175 enable_0/and_6/w_26_9# Gnd 0.82fF
C2176 enable_0/and_6/w_n43_8# Gnd 0.82fF
C2177 enable_0/and_7/a_n26_14# Gnd 0.05fF
C2178 enable_0/en Gnd 3.37fF
C2179 enable_0/and_7/w_26_9# Gnd 0.82fF
C2180 enable_0/and_7/w_n43_8# Gnd 0.82fF
C2181 b1out_0 Gnd 2.82fF
C2182 enable_0/and_5/a_n26_14# Gnd 0.05fF
C2183 enable_0/and_5/w_26_9# Gnd 0.82fF
C2184 enable_0/and_5/w_n43_8# Gnd 0.82fF

.tran 0.1n 200n
.control
run

plot v(a0) v(a1)+2 v(a2)+4 v(a3)+6
plot v(b0) v(b1)+2 v(b2)+4 v(b3)+6
plot v(a0out_2) v(a1out_2)+2 v(a2out_2)+4 v(a3out_2)+6
plot v(b0out_2) v(b1out_2)+2 v(b2out_2)+4 v(b3out_2)+6
* plot v(s0_add) v(s1_add)+2 v(s2_add)+4 v(s3_add)+6 v(fc_add)+8
* plot v(s0_sub) v(s1_sub)+2 v(s2_sub)+4 v(s3_sub)+6 v(fc_sub)+8
* plot v(out0) v(out1)+2 v(out2)+4 v(out3)+6
plot v(equal) v(agb)+2 v(bga)+4

.endc

.end
