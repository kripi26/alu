* SPICE3 file created from 4input_OR.ext - technology: scmos
.include TSMC_180nm.txt
.param SUPPLY = 1.8
.param LAMBDA = 0.09u
.param width_P = 8*LAMBDA
.param width_N = 4*LAMBDA
.global gnd vdd
.option scale=0.09u

Vdd vdd gnd 1.8
va a gnd DC 0
vb b gnd DC 1.8
vc c gnd DC 0
vd d gnd DC 0


M1000 out y vdd NOT_0/vdd CMOSP w=8 l=4
+  ad=101 pd=42 as=199 ps=84
M1001 out y gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=1499 ps=344
M1002 vdd a vdd vdd CMOSP w=14 l=5
+  ad=0 pd=0 as=126 ps=46
M1003 y a gnd Gnd CMOSN w=16 l=7
+  ad=704 pd=216 as=0 ps=0
M1004 vdd c vdd vdd CMOSP w=14 l=5
+  ad=210 pd=58 as=196 ps=56
M1005 y d gnd Gnd CMOSN w=16 l=7
+  ad=0 pd=0 as=0 ps=0
M1006 y b gnd Gnd CMOSN w=16 l=7
+  ad=0 pd=0 as=0 ps=0
M1007 vdd b vdd vdd CMOSP w=14 l=5
+  ad=0 pd=0 as=0 ps=0
M1008 vdd d y vdd CMOSP w=14 l=5
+  ad=0 pd=0 as=238 ps=62
M1009 y c gnd Gnd CMOSN w=16 l=7
+  ad=0 pd=0 as=0 ps=0
C0 a Gnd 4.35fF

.tran 0.1n 500n

.measure tran trise
+ TRIG v(a) VAL = 0.9 RISE = 1
+ TARG v(out) VAL = 0.9 FALL = 1

.measure tran tfall
+ TRIG v(a) VAL = 0.9 FALL = 1
+ TARG v(out) VAL = 0.9 RISE = 1

.measure tran tpd param = '(trise + tfall)/2' goal = 0

.control
run
plot  v(a) v(b)+2 v(c)+4 v(d)+6 v(out)+8
.endc

.end
