magic
tech scmos
timestamp 1700576303
<< polysilicon >>
rect -17 146 4 151
rect -20 88 55 93
rect 2680 -38 2705 -34
rect 4065 -90 4085 -84
rect 1337 -103 1360 -98
rect 2645 -100 2755 -94
rect 4048 -151 4135 -144
rect 1268 -162 1411 -158
<< polycontact >>
rect -21 146 -17 151
rect -25 88 -20 93
rect 2676 -38 2680 -34
rect 4060 -90 4065 -84
rect 1332 -103 1337 -98
rect 2636 -100 2645 -94
rect 4035 -151 4048 -144
rect 1262 -162 1268 -158
<< metal1 >>
rect 47 631 688 639
rect 47 194 52 631
rect 680 553 688 631
rect 4110 618 4774 619
rect 2730 604 3278 615
rect 3744 606 4111 618
rect 4116 606 4775 618
rect 2730 564 2736 604
rect 4768 579 4775 606
rect 1058 551 1387 561
rect 1392 551 1841 561
rect 2307 555 2736 564
rect 382 468 419 472
rect 1621 468 1668 475
rect 604 248 756 254
rect 294 156 299 247
rect 1177 182 1512 188
rect 146 152 299 156
rect -40 146 -21 151
rect -65 88 -25 93
rect -65 -98 -57 88
rect -42 56 -37 88
rect 28 76 32 80
rect 28 74 33 76
rect 13 64 17 66
rect 334 56 595 57
rect -42 49 595 56
rect 334 48 595 49
rect 1387 -54 1392 148
rect 1387 -58 1391 -54
rect 1600 -95 1612 400
rect 2731 308 2736 555
rect 3043 516 3096 526
rect 4552 492 4588 498
rect 5203 488 5206 495
rect 1904 256 2000 257
rect 1904 252 2005 256
rect 2382 184 2886 194
rect 2731 7 2736 151
rect 2957 -25 2971 450
rect 3300 319 3415 333
rect 3402 308 3415 319
rect 3402 303 3443 308
rect 3861 236 4432 242
rect 2659 -38 2676 -34
rect 2847 -35 2971 -25
rect 4111 -43 4116 4
rect 4497 -79 4520 417
rect 4815 274 4925 280
rect 5351 208 5388 214
rect 4032 -90 4060 -84
rect 4227 -87 4520 -79
rect -65 -103 1268 -98
rect 1309 -103 1332 -98
rect 1502 -102 1612 -95
rect 1600 -103 1612 -102
rect 1262 -138 1268 -103
rect 1230 -146 1268 -138
rect 1230 -218 1238 -146
rect 1262 -158 1268 -146
rect 2636 -158 2645 -100
rect 2729 -113 2735 -107
rect 4035 -158 4048 -151
rect 1383 -178 1391 -172
rect 2636 -174 4048 -158
rect 4108 -163 4115 -157
rect 2636 -218 2645 -174
rect 1230 -228 2645 -218
<< m2contact >>
rect 4111 606 4116 618
rect 1387 551 1392 561
rect 1025 462 1034 469
rect 2274 465 2283 472
rect 1600 400 1612 413
rect 1713 400 1722 413
rect 294 247 299 254
rect 464 247 473 254
rect 595 248 604 254
rect 1512 182 1521 188
rect 1387 148 1392 157
rect 28 69 33 74
rect 595 48 604 58
rect 3713 516 3721 523
rect 5206 488 5213 495
rect 2731 302 2736 308
rect 2957 450 2971 464
rect 3151 450 3160 464
rect 1896 252 1904 257
rect 2886 184 2896 194
rect 2731 151 2736 164
rect 4497 417 4520 436
rect 4633 417 4642 436
rect 3280 319 3300 333
rect 4432 236 4437 242
rect 4111 4 4116 10
rect 4807 274 4815 280
rect 2729 -118 2735 -113
rect 1383 -183 1391 -178
rect 4108 -168 4115 -163
<< metal2 >>
rect 1034 462 1218 469
rect 299 247 464 254
rect 13 69 28 74
rect 13 11 18 69
rect 595 58 604 248
rect 1387 157 1392 551
rect 3721 516 3826 523
rect 2283 465 2384 472
rect 2971 450 3151 464
rect 1612 400 1713 413
rect 3050 319 3280 333
rect 1896 188 1904 252
rect 1521 182 1904 188
rect 2731 164 2736 302
rect 3051 194 3064 319
rect 2896 185 3064 194
rect 2896 184 3062 185
rect 761 11 769 73
rect 13 4 769 11
rect 809 -302 831 70
rect 1383 -302 1391 -183
rect 809 -304 1391 -302
rect 2048 -301 2079 71
rect 2729 -301 2735 -118
rect 3555 -301 3573 128
rect 4111 10 4116 606
rect 5213 488 5255 495
rect 4520 417 4633 436
rect 4807 242 4815 274
rect 4437 236 4815 242
rect 4108 -301 4115 -168
rect 2048 -302 4115 -301
rect 4998 -302 5010 99
rect 2048 -304 5010 -302
rect 809 -319 5010 -304
rect 1379 -320 5010 -319
rect 1379 -321 5009 -320
use fulladder  fulladder_3
timestamp 1700494352
transform 1 0 4742 0 1 391
box -164 -302 611 196
use XOR  XOR_3
timestamp 1699220400
transform 1 0 4122 0 1 -88
box -56 -86 137 64
use fulladder  fulladder_2
timestamp 1700494352
transform 1 0 3260 0 1 419
box -164 -302 611 196
use XOR  XOR_2
timestamp 1699220400
transform 1 0 2742 0 1 -38
box -56 -86 137 64
use fulladder  fulladder_1
timestamp 1700494352
transform 1 0 1822 0 1 368
box -164 -302 611 196
use XOR  XOR_1
timestamp 1699220400
transform 1 0 1397 0 1 -103
box -56 -86 137 64
use fulladder  fulladder_0
timestamp 1700494352
transform 1 0 573 0 1 365
box -164 -302 611 196
use XOR  XOR_0
timestamp 1699220400
transform 1 0 41 0 1 149
box -56 -86 137 64
<< labels >>
rlabel metal1 -28 148 -27 149 1 b0
rlabel metal1 -30 90 -29 91 1 M
rlabel metal1 393 469 394 470 1 a0
rlabel metal1 1204 184 1205 185 1 c1
rlabel metal1 1624 471 1625 472 1 a1
rlabel metal2 2365 467 2366 468 1 s1
rlabel metal1 2485 187 2487 189 1 c2
rlabel metal1 2670 -37 2671 -36 1 b2
rlabel metal1 3060 519 3061 520 1 a2
rlabel metal2 3799 518 3800 519 1 s2
rlabel metal1 3890 238 3891 240 1 c3
rlabel metal1 4048 -88 4051 -86 1 b3
rlabel metal1 4564 494 4565 495 1 a3
rlabel metal2 5247 490 5248 492 1 s3
rlabel metal1 5377 211 5378 212 1 c4
rlabel metal1 354 633 356 636 5 vdd
rlabel metal2 475 7 477 8 1 gnd
rlabel metal1 197 153 198 154 1 b0xorM
rlabel metal2 1205 465 1205 465 1 s0
rlabel metal1 1317 -100 1317 -100 1 b1
rlabel space 757 469 757 469 1 a0xorb0
rlabel space 916 135 916 135 1 ab
<< end >>
