.include TSMC_180nm.txt
.include "AND.sub"
.include "NOT.sub"

.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd node_x gnd 'SUPPLY'

V_in_a node_a gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 40ns)
V_in_b node_b gnd PULSE(0 1.8 0ns 100ps 100ps 50ns 70ns)

X1 node_a node_c node_x gnd NOT
X2 node_b node_d node_x gnd NOT     

* node_b - S1
* node_a - S0

X3 node_c node_d node_out0 node_x gnd AND
X4 node_a node_d node_out1 node_x gnd AND
X5 node_b node_c node_out2 node_x gnd AND
X6 node_a node_b node_out3 node_x gnd AND

C1 node_out0 gnd 100f
C2 node_out1 gnd 100f
C3 node_out2 gnd 100f
C4 node_out3 gnd 100f



.tran 1n 800n


.control
run
set color0 = rgb:f/f/e
set color1 = white
plot v(node_a) v(node_b)+2 v(node_out3)+4
plot v(node_a) v(node_b)+2 v(node_out2)+4
plot v(node_a) v(node_b)+2 v(node_out1)+4
plot v(node_a) v(node_b)+2 v(node_out0)+4
* hardcopy image.ps v(node_a) v(node_b)+2 v(node_out)+4
.end
.endc

