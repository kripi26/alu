magic
tech scmos
timestamp 1700972767
<< polysilicon >>
rect 3 88 12 92
rect 0 -13 12 -9
rect 0 -114 12 -110
rect 0 -212 12 -208
<< polycontact >>
rect -1 88 3 92
rect 21 75 25 79
rect -5 -13 0 -9
rect 21 -25 25 -21
rect -5 -114 0 -110
rect 21 -124 25 -120
rect -5 -212 0 -208
rect 21 -223 25 -219
<< metal1 >>
rect -43 117 5 122
rect -43 22 -37 117
rect -20 88 -1 92
rect 97 84 120 88
rect -16 75 21 79
rect 112 48 160 55
rect -43 16 3 22
rect -43 -77 -37 16
rect -23 -13 -5 -9
rect 97 -18 120 -14
rect -16 -25 21 -21
rect 154 -45 160 48
rect 112 -52 160 -45
rect -43 -83 6 -77
rect -43 -176 -37 -83
rect -23 -114 -5 -110
rect 97 -117 120 -113
rect -16 -124 21 -120
rect 154 -144 160 -52
rect 111 -151 160 -144
rect -43 -181 4 -176
rect -21 -212 -5 -208
rect 97 -215 120 -211
rect -16 -223 21 -219
rect 154 -243 160 -151
rect 111 -250 160 -243
use and  and_3
timestamp 1699973769
transform 1 0 38 0 1 -212
box -43 -38 74 36
use and  and_2
timestamp 1699973769
transform 1 0 38 0 1 -113
box -43 -38 74 36
use and  and_1
timestamp 1699973769
transform 1 0 38 0 1 -14
box -43 -38 74 36
use and  and_0
timestamp 1699973769
transform 1 0 38 0 1 86
box -43 -38 74 36
<< labels >>
rlabel metal1 -8 91 -8 91 1 a0
rlabel metal1 0 77 0 77 1 b0
rlabel metal1 -9 -12 -9 -12 1 a1
rlabel metal1 2 -24 2 -24 1 b1
rlabel metal1 -9 -112 -9 -112 1 a2
rlabel metal1 4 -122 4 -122 1 b2
rlabel metal1 -10 -211 -10 -211 1 a3
rlabel metal1 0 -220 0 -220 1 b3
rlabel metal1 117 86 117 86 7 y0
rlabel metal1 115 -16 115 -16 7 y1
rlabel metal1 115 -116 115 -116 7 y2
rlabel metal1 114 -214 114 -214 1 y3
rlabel metal1 -19 119 -19 119 5 vdd
rlabel metal1 144 -246 144 -246 1 gnd
<< end >>
