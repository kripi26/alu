magic
tech scmos
timestamp 1701544513
<< metal1 >>
rect 1495 2284 1515 2285
rect 753 2261 1515 2284
rect 849 2155 878 2156
rect -50 2140 878 2155
rect -50 315 -44 2140
rect 692 2139 713 2140
rect 106 2044 586 2054
rect 607 2044 642 2054
rect 106 417 110 2044
rect 636 1947 642 2044
rect 775 1914 783 1918
rect 645 1906 655 1910
rect 766 1781 844 1785
rect 641 1775 644 1780
rect 767 1674 836 1678
rect 639 1667 645 1672
rect 767 1565 827 1569
rect 639 1558 643 1564
rect 780 1447 781 1449
rect 767 1443 781 1447
rect 640 1435 645 1441
rect 767 1341 781 1345
rect 638 1333 645 1338
rect 752 1242 781 1246
rect 638 1240 645 1241
rect 638 1236 656 1240
rect 780 1146 781 1147
rect 754 1142 781 1146
rect 612 1141 640 1142
rect 612 1137 641 1141
rect 775 990 816 994
rect 641 982 645 987
rect 766 857 808 861
rect 639 851 644 856
rect 767 750 800 754
rect 639 743 645 748
rect 767 641 794 645
rect 638 634 643 639
rect 766 519 781 523
rect 639 511 644 517
rect 765 417 781 423
rect 640 409 645 414
rect -50 310 -15 315
rect 637 312 644 318
rect 611 213 642 218
rect 632 43 637 167
rect 791 99 794 641
rect 797 109 800 750
rect 803 200 808 857
rect 812 685 816 990
rect 822 967 827 1565
rect 831 1398 836 1674
rect 840 1413 844 1781
rect 849 1570 878 2140
rect 1495 2071 1515 2261
rect 5852 1931 5962 1937
rect 2718 1907 3031 1914
rect 5852 1643 5859 1931
rect 6795 1647 6803 1653
rect 849 1532 877 1570
rect 849 1527 1355 1532
rect 2709 1413 2718 1501
rect 840 1406 1245 1413
rect 1658 1406 2718 1413
rect 3985 1401 4068 1405
rect 831 1392 1187 1398
rect 1180 1084 1187 1392
rect 2213 1344 2250 1352
rect 1344 1211 1352 1341
rect 2096 1242 2620 1247
rect 3985 1247 3991 1401
rect 5373 1349 5443 1355
rect 2777 1241 3991 1247
rect 3924 1107 3933 1147
rect 1180 1078 3924 1084
rect 5362 1066 5373 1233
rect 5852 967 5859 1293
rect 822 963 5859 967
rect 5881 705 5994 711
rect 2919 681 3061 688
rect 812 679 816 680
rect 2919 579 2936 681
rect 2681 568 2936 579
rect 5881 354 5889 705
rect 6826 421 6834 427
rect 2180 190 2352 200
rect 2195 161 2758 169
rect 2748 109 2758 161
rect 797 105 1345 109
rect 791 95 1321 99
rect 801 38 1267 42
rect 279 -1817 286 3
rect 360 -941 367 34
rect 668 30 671 35
rect 791 -95 1243 -88
rect 668 -101 671 -96
rect 792 -202 1222 -195
rect 667 -209 671 -204
rect 788 -311 1203 -301
rect 666 -318 668 -313
rect 787 -433 851 -425
rect 665 -441 671 -435
rect 787 -535 1127 -526
rect 663 -543 671 -537
rect 778 -634 993 -622
rect 663 -640 670 -634
rect 780 -734 1101 -728
rect 629 -739 668 -734
rect 360 -945 637 -941
rect 1072 -944 1087 -943
rect 798 -950 1088 -944
rect 665 -958 671 -953
rect 786 -1083 1065 -1075
rect 667 -1089 672 -1084
rect 788 -1190 1046 -1183
rect 668 -1197 671 -1192
rect 787 -1299 1032 -1294
rect 666 -1306 669 -1301
rect 788 -1421 1016 -1415
rect 666 -1429 671 -1423
rect 787 -1523 1003 -1515
rect 663 -1531 671 -1525
rect 774 -1622 991 -1615
rect 664 -1628 670 -1623
rect 632 -1727 669 -1721
rect 778 -1722 968 -1715
rect 711 -1817 721 -1748
rect 279 -1826 721 -1817
rect 958 -5412 968 -1722
rect 982 -5313 991 -1622
rect 996 -5215 1003 -1523
rect 1009 -5114 1015 -1421
rect 1027 -5401 1032 -1299
rect 1040 -5241 1046 -1190
rect 1055 -5180 1065 -1083
rect 1072 -5101 1087 -950
rect 1191 -2336 1203 -311
rect 1213 -2574 1222 -202
rect 1230 -291 1243 -95
rect 1254 -173 1267 38
rect 1230 -2812 1244 -291
rect 1253 -2943 1268 -173
rect 1317 -249 1321 95
rect 1337 -216 1345 105
rect 3991 -216 4000 -47
rect 1337 -224 4000 -216
rect 5881 -249 5889 46
rect 1317 -254 5889 -249
rect 3969 -1379 3977 -1376
rect 3420 -2755 3443 -2752
rect 1253 -3087 1269 -2943
rect 1253 -3095 2090 -3087
rect 3949 -4080 3965 -4077
rect 2388 -5080 2394 -4994
rect 2463 -5111 2467 -5107
rect 2497 -5148 2503 -4548
rect 1054 -5198 1065 -5180
rect 2461 -5213 2469 -5209
rect 1039 -5303 1046 -5241
rect 2463 -5312 2467 -5308
rect 2463 -5410 2467 -5406
rect 958 -5419 2332 -5412
<< m2contact >>
rect 713 2261 753 2284
rect 586 2044 607 2054
rect 783 1914 788 1919
rect 640 1906 645 1911
rect 636 1775 641 1780
rect 634 1667 639 1672
rect 634 1558 639 1564
rect 781 1443 788 1449
rect 634 1435 640 1441
rect 781 1341 787 1347
rect 632 1333 638 1338
rect 781 1242 787 1247
rect 633 1236 638 1241
rect 605 1187 610 1201
rect 781 1142 786 1147
rect 607 1137 612 1142
rect 754 1110 759 1117
rect 636 982 641 987
rect 754 955 759 962
rect 634 851 639 856
rect 633 743 639 748
rect 632 634 638 639
rect 781 519 786 524
rect 634 511 639 517
rect 781 417 787 423
rect 634 409 640 415
rect 279 384 286 390
rect 748 318 753 323
rect 632 312 637 318
rect 291 264 299 269
rect 605 264 610 269
rect 750 218 755 223
rect 606 213 611 218
rect 749 186 756 193
rect 324 167 330 173
rect 632 167 637 173
rect 4452 1955 4470 1965
rect 1791 1907 1796 1912
rect 2709 1907 2718 1914
rect 5852 1637 5859 1643
rect 1364 1585 1370 1591
rect 2709 1501 2719 1510
rect 1245 1406 1253 1413
rect 1650 1406 1658 1413
rect 2203 1344 2213 1352
rect 2250 1344 2260 1352
rect 2718 1336 2724 1341
rect 2086 1242 2096 1248
rect 2620 1242 2626 1248
rect 5362 1349 5373 1355
rect 2770 1241 2777 1247
rect 5852 1293 5859 1298
rect 1344 1203 1352 1211
rect 5362 1233 5373 1246
rect 3924 1147 3933 1155
rect 3924 1101 3933 1107
rect 3924 1078 3933 1084
rect 5362 1056 5373 1066
rect 1491 844 1496 852
rect 4483 728 4494 739
rect 812 680 817 685
rect 1822 680 1838 685
rect 2671 568 2681 579
rect 1400 359 1405 368
rect 5881 346 5889 354
rect 1375 297 1383 306
rect 803 190 808 200
rect 2170 190 2180 200
rect 2352 190 2362 201
rect 4099 175 4107 183
rect 2184 161 2195 169
rect 5472 123 5477 131
rect 663 30 668 35
rect 776 3 784 10
rect 662 -101 668 -96
rect 661 -209 667 -204
rect 660 -318 666 -313
rect 851 -433 860 -425
rect 659 -441 665 -435
rect 1127 -535 1143 -526
rect 658 -543 663 -537
rect 993 -634 1005 -621
rect 658 -640 663 -634
rect 623 -739 629 -734
rect 1101 -738 1114 -728
rect 779 -766 784 -759
rect 660 -958 665 -953
rect 779 -985 784 -978
rect 661 -1089 667 -1084
rect 663 -1197 668 -1192
rect 660 -1306 666 -1301
rect 660 -1429 666 -1423
rect 658 -1531 663 -1525
rect 659 -1628 664 -1623
rect 627 -1727 632 -1721
rect 1009 -5122 1015 -5114
rect 996 -5220 1003 -5215
rect 982 -5320 991 -5313
rect 1190 -2351 1203 -2336
rect 1213 -2582 1222 -2574
rect 1230 -2823 1244 -2812
rect 5881 46 5889 54
rect 3991 -47 4000 -35
rect 2425 -892 2432 -885
rect 2388 -4994 2394 -4987
rect 1072 -5108 1087 -5101
rect 2323 -5107 2328 -5101
rect 2327 -5120 2333 -5114
rect 1054 -5208 1066 -5198
rect 2320 -5208 2329 -5200
rect 2327 -5220 2336 -5215
rect 1039 -5308 1046 -5303
rect 2320 -5308 2328 -5303
rect 2327 -5320 2332 -5313
rect 1027 -5407 1032 -5401
rect 2322 -5407 2327 -5401
<< metal2 >>
rect 586 2284 607 2285
rect 586 2261 713 2284
rect 586 2054 607 2261
rect 3923 1955 4452 1965
rect 5229 1955 5250 1962
rect 3923 1954 4470 1955
rect 788 1914 1750 1919
rect 1746 1911 1750 1914
rect 2709 1914 2718 1915
rect 631 1906 640 1911
rect 1746 1907 1791 1911
rect 2612 1900 2649 1908
rect 634 1775 636 1780
rect 631 1667 634 1672
rect 1156 1591 1165 1592
rect 1156 1585 1364 1591
rect 632 1558 634 1564
rect 1156 1449 1165 1585
rect 2709 1510 2718 1907
rect 3788 1904 3809 1911
rect 788 1443 1165 1449
rect 633 1435 634 1441
rect 1253 1406 1650 1413
rect 787 1344 2203 1347
rect 787 1341 2213 1344
rect 2260 1344 2724 1347
rect 2250 1341 2724 1344
rect 631 1333 632 1338
rect 787 1242 2086 1247
rect 2626 1242 2770 1247
rect 2620 1241 2770 1242
rect 631 1236 633 1241
rect 343 1187 605 1201
rect 344 390 355 1187
rect 583 1137 607 1142
rect 617 1094 622 1184
rect 786 1142 982 1147
rect 617 1023 622 1087
rect 754 1046 759 1110
rect 977 1066 982 1142
rect 1344 1112 1352 1203
rect 3924 1155 3933 1954
rect 6661 1927 6676 1934
rect 5362 1246 5373 1349
rect 5852 1298 5859 1637
rect 3924 1084 3933 1101
rect 977 1056 5362 1066
rect 754 1041 2361 1046
rect 406 982 590 987
rect 634 982 636 987
rect 754 962 759 1041
rect 908 897 1496 906
rect 421 851 595 856
rect 631 851 634 856
rect 1491 852 1496 897
rect 442 743 592 748
rect 632 743 633 748
rect 3991 728 4483 739
rect 5266 729 5279 736
rect 817 680 1822 685
rect 2651 675 2667 682
rect 3824 678 3833 685
rect 458 634 593 639
rect 631 634 632 639
rect 786 519 1312 524
rect 482 511 593 517
rect 631 511 634 517
rect 493 409 587 415
rect 632 409 634 415
rect 286 384 355 390
rect 753 318 756 323
rect 547 312 594 318
rect 631 312 632 318
rect 299 264 605 269
rect 583 213 606 218
rect -30 189 4 194
rect 617 181 622 263
rect 755 218 757 223
rect 617 178 648 181
rect 330 167 632 173
rect 643 71 648 178
rect 749 118 756 186
rect 781 169 787 417
rect 1305 368 1312 519
rect 1305 359 1400 368
rect 1344 306 1352 334
rect 1344 297 1375 306
rect 808 190 2170 200
rect 2671 200 2681 568
rect 2362 190 2681 200
rect 781 161 2184 169
rect 749 109 784 118
rect 776 62 784 109
rect 776 52 2271 62
rect 406 30 597 35
rect 660 30 663 35
rect 776 10 784 52
rect 776 2 784 3
rect 3991 -35 4000 728
rect 6694 701 6736 708
rect 4027 175 4099 183
rect 5399 123 5472 131
rect 5881 54 5889 346
rect 421 -101 591 -96
rect 658 -101 662 -96
rect 441 -208 596 -204
rect 433 -209 596 -208
rect 659 -209 661 -204
rect 458 -318 593 -313
rect 658 -318 660 -313
rect 860 -433 1313 -425
rect 482 -441 611 -435
rect 657 -441 659 -435
rect 1143 -535 1184 -526
rect 493 -542 587 -537
rect 488 -543 587 -542
rect 657 -543 658 -537
rect 1176 -597 1184 -535
rect 1005 -634 1152 -621
rect 547 -640 605 -634
rect 657 -640 658 -634
rect 583 -739 623 -734
rect 643 -824 648 -692
rect 643 -917 648 -835
rect 779 -759 784 -758
rect 779 -886 784 -766
rect 406 -958 602 -953
rect 658 -958 660 -953
rect 779 -978 784 -892
rect 1104 -924 1114 -738
rect 1103 -1004 1114 -924
rect 1143 -781 1152 -634
rect 1175 -701 1184 -597
rect 421 -1089 598 -1084
rect 659 -1089 661 -1084
rect 442 -1197 608 -1192
rect 661 -1197 663 -1192
rect 458 -1306 617 -1301
rect 659 -1306 660 -1301
rect 482 -1429 590 -1423
rect 658 -1429 660 -1423
rect 493 -1531 596 -1525
rect 657 -1531 658 -1525
rect 1103 -1550 1115 -1004
rect 1143 -1399 1153 -781
rect 1174 -984 1184 -701
rect 1304 -823 1313 -433
rect 1304 -856 1314 -823
rect 1304 -867 2139 -856
rect 2360 -892 2425 -886
rect 1174 -1135 1183 -984
rect 1174 -1156 1970 -1135
rect 1144 -1454 1153 -1399
rect 547 -1628 608 -1623
rect 658 -1628 659 -1623
rect 583 -1727 627 -1721
rect 1104 -1722 1115 -1550
rect 1203 -2351 1996 -2336
rect 1222 -2582 2053 -2574
rect 2266 -2582 2287 -2572
rect 1761 -2812 2056 -2811
rect 1244 -2823 2056 -2812
rect 2388 -4987 2394 -4908
rect 1087 -5107 2323 -5101
rect 1015 -5120 2327 -5114
rect 1015 -5122 2331 -5120
rect 1066 -5208 2320 -5200
rect 1003 -5220 2327 -5215
rect 1046 -5308 2320 -5303
rect 991 -5320 2327 -5313
rect 1032 -5407 2322 -5401
<< m3contact >>
rect 626 1906 631 1911
rect 629 1775 634 1780
rect 626 1667 631 1672
rect 626 1558 632 1564
rect 628 1435 633 1441
rect 626 1333 631 1338
rect 626 1236 631 1241
rect 577 1137 583 1142
rect 617 1087 622 1094
rect 2361 1120 2369 1137
rect 1344 1104 1352 1112
rect 2361 1041 2369 1046
rect 401 982 406 987
rect 590 982 595 987
rect 629 982 634 987
rect 903 897 908 906
rect 415 851 421 856
rect 595 851 600 856
rect 626 851 631 856
rect 433 743 442 748
rect 592 743 597 748
rect 626 743 632 748
rect 452 634 458 639
rect 593 634 599 639
rect 626 634 631 639
rect 474 511 482 517
rect 593 511 598 517
rect 626 511 631 517
rect 488 409 493 415
rect 587 409 592 415
rect 626 409 632 415
rect 756 318 761 323
rect 541 312 547 318
rect 594 312 599 318
rect 626 312 631 318
rect 577 213 583 218
rect 757 218 762 223
rect 1344 334 1352 346
rect 401 30 406 35
rect 597 30 602 35
rect 655 30 660 35
rect 4016 175 4027 183
rect 5388 123 5399 131
rect 415 -101 421 -96
rect 591 -101 597 -96
rect 653 -101 658 -96
rect 432 -208 441 -203
rect 596 -209 601 -204
rect 654 -209 659 -204
rect 452 -318 458 -313
rect 593 -318 599 -313
rect 652 -318 658 -313
rect 474 -441 482 -435
rect 611 -441 618 -435
rect 652 -441 657 -435
rect 488 -542 493 -537
rect 587 -543 592 -537
rect 652 -543 657 -537
rect 541 -640 547 -634
rect 605 -640 610 -634
rect 652 -640 657 -634
rect 577 -739 583 -734
rect 643 -835 648 -824
rect 778 -892 784 -886
rect 401 -958 406 -953
rect 602 -958 608 -953
rect 653 -958 658 -953
rect 415 -1089 421 -1084
rect 598 -1089 604 -1084
rect 653 -1089 659 -1084
rect 433 -1197 442 -1192
rect 608 -1197 613 -1192
rect 656 -1197 661 -1192
rect 452 -1306 458 -1301
rect 617 -1306 622 -1301
rect 653 -1306 659 -1301
rect 474 -1429 482 -1423
rect 590 -1429 595 -1423
rect 652 -1429 658 -1423
rect 488 -1531 493 -1525
rect 596 -1531 601 -1525
rect 652 -1531 657 -1525
rect 2354 -892 2360 -886
rect 1970 -1156 1986 -1132
rect 2169 -1156 2181 -1140
rect 1144 -1461 1153 -1454
rect 2230 -1467 2243 -1461
rect 541 -1628 547 -1623
rect 608 -1628 614 -1623
rect 652 -1628 658 -1623
rect 577 -1727 583 -1721
rect 1104 -1737 1115 -1722
rect 2279 -1737 2286 -1723
rect 1996 -2351 2005 -2336
rect 2053 -2582 2063 -2574
rect 2259 -2582 2266 -2572
rect 2056 -2823 2068 -2811
rect 2197 -2823 2207 -2811
rect 2411 -4107 2416 -4100
rect 2388 -4908 2394 -4901
<< metal3 >>
rect 401 1906 626 1911
rect 401 987 406 1906
rect 401 35 406 982
rect 401 -953 406 30
rect 415 1775 629 1780
rect 415 856 421 1775
rect 415 -96 421 851
rect 415 -1084 421 -101
rect 433 1667 626 1672
rect 433 748 442 1667
rect 433 -203 442 743
rect 441 -208 442 -203
rect 433 -1192 442 -208
rect 452 1558 626 1564
rect 452 639 458 1558
rect 452 -313 458 634
rect 452 -1301 458 -318
rect 474 1435 628 1441
rect 474 517 482 1435
rect 474 -435 482 511
rect 474 -1423 482 -441
rect 488 1333 626 1338
rect 488 415 493 1333
rect 488 -537 493 409
rect 488 -1525 493 -542
rect 541 1236 626 1241
rect 541 318 547 1236
rect 541 -634 547 312
rect 541 -1623 547 -640
rect 577 218 583 1137
rect 903 1094 908 1095
rect 622 1087 908 1094
rect 595 982 629 987
rect 903 906 908 1087
rect 600 851 626 856
rect 597 743 626 748
rect 599 634 626 639
rect 598 511 626 517
rect 592 409 626 415
rect 1344 346 1352 1104
rect 2361 1046 2369 1120
rect 761 318 1320 323
rect 599 312 626 318
rect 762 218 1281 223
rect 577 -734 583 213
rect 1274 92 1281 218
rect 1312 131 1320 318
rect 1312 124 2582 131
rect 1274 86 2103 92
rect 602 30 655 35
rect 597 -101 653 -96
rect 2097 -111 2103 86
rect 2572 -63 2582 124
rect 4016 -63 4027 175
rect 2572 -70 4027 -63
rect 5388 -111 5399 123
rect 2097 -117 5399 -111
rect 601 -209 654 -204
rect 599 -318 652 -313
rect 618 -441 652 -435
rect 1403 -457 1417 -455
rect 1402 -479 2769 -457
rect 592 -543 652 -537
rect 610 -640 652 -634
rect 577 -1721 583 -739
rect 1403 -824 1417 -479
rect 648 -835 1417 -824
rect 784 -892 2354 -886
rect 608 -958 653 -953
rect 604 -1089 653 -1084
rect 1986 -1140 2181 -1132
rect 1986 -1156 2169 -1140
rect 613 -1197 656 -1192
rect 622 -1306 653 -1301
rect 595 -1429 652 -1423
rect 1960 -1454 2243 -1453
rect 1153 -1461 2243 -1454
rect 601 -1531 652 -1525
rect 614 -1628 652 -1623
rect 1115 -1737 2279 -1723
rect 2063 -2582 2259 -2574
rect 2068 -2823 2197 -2811
rect 2388 -4107 2411 -4100
rect 2388 -4901 2394 -4107
use comparator  comparator_0
timestamp 1701538741
transform 1 0 2474 0 1 -2442
box -478 -2141 1498 1985
use enable  enable_3
timestamp 1701496846
transform 1 0 703 0 1 -996
box -71 -758 100 85
use enable  enable_2
timestamp 1701496846
transform 1 0 703 0 1 -8
box -71 -758 100 85
use enable  enable_1
timestamp 1701496846
transform 1 0 677 0 1 944
box -71 -758 100 85
use enable  enable_0
timestamp 1701496846
transform 1 0 677 0 1 1868
box -71 -758 100 85
use 4bitadder  4bitadder_0
timestamp 1700576303
transform 1 0 1409 0 1 1439
box -65 -321 5388 639
use decoder  decoder_0
timestamp 1700447719
transform 1 0 69 0 1 230
box -93 -233 302 193
use 4bitadder  4bitadder_1
timestamp 1700576303
transform 1 0 1440 0 1 213
box -65 -321 5388 639
use AND_Block  AND_Block_0
timestamp 1700972767
transform 1 0 2343 0 1 -5195
box -43 -250 160 122
<< labels >>
rlabel metal1 -30 312 -30 312 1 s0
rlabel metal2 -25 192 -25 192 1 s1
rlabel metal3 614 1560 614 1560 1 a3
rlabel metal1 621 1139 621 1139 1 b3
rlabel metal1 778 1144 778 1144 1 b3out_0
rlabel metal1 779 1244 779 1244 1 b2out_0
rlabel metal1 779 1343 779 1343 1 b1out_0
rlabel metal1 779 1445 779 1445 1 b0out_0
rlabel metal1 779 1567 779 1567 1 a3out_0
rlabel metal1 779 1783 779 1783 1 a1out_0
rlabel metal1 778 1916 778 1916 1 a0out_0
rlabel metal2 636 1908 636 1908 1 a0
rlabel metal1 641 1239 641 1239 1 b2
rlabel metal1 642 1335 642 1335 1 b1
rlabel metal1 642 1437 642 1437 1 b0
rlabel metal1 641 1669 641 1669 1 a2
rlabel metal1 643 1778 643 1778 1 a1
rlabel metal1 575 2047 575 2047 1 vdd
rlabel metal1 600 -1823 600 -1823 1 gnd
rlabel metal1 2463 -5111 2467 -5107 1 out0
rlabel metal1 2463 -5312 2467 -5308 1 out2
rlabel metal1 2463 -5410 2467 -5406 1 out3
rlabel metal1 2463 -5213 2469 -5209 1 out1
rlabel metal1 3974 -1377 3974 -1377 1 agb
rlabel metal1 3439 -2753 3439 -2753 1 equal
rlabel metal1 3963 -4078 3963 -4078 1 bga
rlabel metal2 2662 679 2662 679 1 s0_sub
rlabel metal2 3828 682 3828 682 1 s1_sub
rlabel metal2 5275 733 5275 733 1 s2_sub
rlabel metal2 6718 705 6719 706 1 s3_sub
rlabel metal2 2642 1906 2642 1906 1 s0_add
rlabel metal2 3804 1907 3804 1907 1 s1_add
rlabel metal2 5237 1959 5237 1959 1 s2_add
rlabel metal2 6672 1931 6672 1931 1 s3_add
rlabel metal1 6799 1650 6799 1650 1 fc_add
rlabel metal1 6829 424 6829 424 7 fc_sub
rlabel metal1 787 1676 787 1676 1 a2out_0
rlabel metal1 811 993 811 993 1 a0_out1
rlabel metal1 804 859 804 859 1 a1out_1
rlabel metal1 797 752 797 752 1 a2out_1
rlabel metal1 790 643 790 643 1 a3out_1
rlabel metal2 788 521 788 521 1 b0out_1
rlabel metal2 784 413 784 413 1 b1out_1
rlabel metal3 766 321 766 321 1 b2out_1
rlabel metal3 765 221 765 221 1 b3out_1
rlabel metal1 1259 38 1259 38 1 a0out_2
rlabel metal1 1234 -92 1234 -92 1 a1out_2
rlabel metal1 1218 -198 1218 -198 1 a2out_2
rlabel metal1 1199 -305 1199 -305 1 a3out_2
rlabel metal1 834 -428 834 -428 1 boout_2
rlabel metal1 825 -529 825 -529 1 b1out_2
rlabel metal1 957 -631 961 -630 1 b2out_2
rlabel metal1 829 -730 829 -730 1 b3out_2
rlabel metal1 863 -946 863 -946 1 a0out_3
rlabel metal1 931 -1079 931 -1079 1 a1out_3
rlabel metal1 935 -1188 935 -1188 1 a2out_3
rlabel metal1 887 -1297 887 -1297 1 a3out_3
rlabel metal1 966 -1418 967 -1417 1 b0out_3
rlabel metal1 911 -1521 912 -1520 1 b1out_3
rlabel metal1 954 -1619 954 -1619 1 b2out_3
rlabel metal1 941 -1719 941 -1719 1 b3out_3
<< end >>
