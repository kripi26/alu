.include TSMC_180nm.txt
.include "decoder.sub"
.include "comparator.sub"
.include "and.sub"
.include "full_adder.sub"
.include "XOR.sub"
.include "enable.sub"
.include "4bitadder.sub"
.include 'AND_block.sub'

.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd node_x gnd 'SUPPLY'

V_in_s0 node_s0 gnd DC 1.8
V_in_s1 node_s1 gnd DC 1.8
V_in_a0 node_a0 gnd DC 0
V_in_a1 node_a1 gnd DC 0
V_in_a2 node_a2 gnd DC 0
V_in_a3 node_a3 gnd DC 1.8
V_in_b0 node_b0 gnd DC 1.8
V_in_b1 node_b1 gnd DC 1.8
V_in_b2 node_b2 gnd DC 1.8
V_in_b3 node_b3 gnd DC 0

X1 node_s0 node_s1 node_out0 node_out1 node_out2 node_out3 node_x gnd decoder

X2 node_a0 node_a1 node_a2 node_a3 node_b0 node_b1 node_b2 node_b3 node_out0 node_a0_out0 node_a1_out0 node_a2_out0 node_a3_out0 node_b0_out0 node_b1_out0 node_b2_out0 node_b3_out0 node_x gnd enable
X3 node_a0 node_a1 node_a2 node_a3 node_b0 node_b1 node_b2 node_b3 node_out1 node_a0_out1 node_a1_out1 node_a2_out1 node_a3_out1 node_b0_out1 node_b1_out1 node_b2_out1 node_b3_out1 node_x gnd enable
X4 node_a0 node_a1 node_a2 node_a3 node_b0 node_b1 node_b2 node_b3 node_out2 node_a0_out2 node_a1_out2 node_a2_out2 node_a3_out2 node_b0_out2 node_b1_out2 node_b2_out2 node_b3_out2 node_x gnd enable
X5 node_a0 node_a1 node_a2 node_a3 node_b0 node_b1 node_b2 node_b3 node_s1 node_a0_out3 node_a1_out3 node_a2_out3 node_a3_out3 node_b0_out3 node_b1_out3 node_b2_out3 node_b3_out3 node_x gnd enable

* 4 bit adder

X6 node_a0_out0 node_a1_out0 node_a2_out0 node_a3_out0 node_b0_out0 node_b1_out0 node_b2_out0 node_b3_out0 node_s0 node_C4_add node_S0_add node_S1_add node_S2_add node_S3_add node_x gnd 4bitadder

* 4 bit subractor
X7 node_a0_out1 node_a1_out1 node_a2_out1 node_a3_out1 node_b0_out1 node_b1_out1 node_b2_out1 node_b3_out1 node_s0 node_C4_sub node_S0_sub node_S1_sub node_S2_sub node_S3_sub node_x gnd 4bitadder


* * comparator
X22 node_a0_out2 node_a1_out2 node_a2_out2 node_a3_out2 node_b0_out2 node_b1_out2 node_b2_out2 node_b3_out2 node_equal node_ab node_ba node_x gnd comparator

* * And block
X8 node_a0_out3 node_a1_out3 node_a2_out3 node_a3_out3 node_b0_out3 node_b1_out3 node_b2_out3 node_b3_out3 node_out0 node_out1 node_out2 node_out3 node_x gnd AND_block


C1 node_C4_add gnd 100f
C2 node_S3_add gnd 100f
C3 node_S2_add gnd 100f
C4 node_S1_add gnd 100f
C5 node_S0_add gnd 100f

.tran 1n 800n


.control
run
set color0 = rgb:f/f/e
set color1 = white
* plot v(node_s0) v(node_s1)+2 
plot v(node_a3) v(node_a2)+2 v(node_a1)+4 v(node_a0)+6
plot v(node_b3) v(node_b2)+2 v(node_b1)+4 v(node_b0)+6
plot v(node_out0) v(node_out1)+2 v(node_out2)+4 v(node_out3)+6
* hardcopy image.ps v(node_a) v(node_b)+2 v(node_out)+4
.end
.endc