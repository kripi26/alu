magic
tech scmos
timestamp 1700474897
<< nwell >>
rect -14 24 11 69
rect 32 -21 57 24
rect 69 -71 94 -26
<< ntransistor >>
rect -9 -97 6 -89
rect -9 -116 6 -108
rect -9 -133 6 -125
<< ptransistor >>
rect -8 45 5 53
rect 38 -1 51 7
rect 75 -50 88 -42
<< ndiffusion >>
rect -9 -85 -5 -78
rect 1 -85 6 -78
rect -9 -89 6 -85
rect -9 -108 6 -97
rect -9 -125 6 -116
rect -9 -138 6 -133
rect -9 -144 -5 -138
rect 2 -144 6 -138
<< pdiffusion >>
rect -8 57 -6 63
rect 1 57 5 63
rect -8 53 5 57
rect -8 38 5 45
rect -8 32 -5 38
rect 1 32 5 38
rect 38 11 41 16
rect 48 11 51 16
rect 38 7 51 11
rect 38 -7 51 -1
rect 44 -13 51 -7
rect 38 -15 51 -13
rect 75 -39 78 -34
rect 85 -39 88 -34
rect 75 -42 88 -39
rect 75 -57 88 -50
rect 81 -63 88 -57
rect 75 -65 88 -63
<< ndcontact >>
rect -5 -85 1 -78
rect -5 -144 2 -138
<< pdcontact >>
rect -6 57 1 63
rect -5 32 1 38
rect 41 11 48 16
rect 38 -13 44 -7
rect 78 -39 85 -34
rect 75 -63 81 -57
<< polysilicon >>
rect -121 45 -8 53
rect 5 45 17 53
rect -121 -125 -114 45
rect -81 -1 38 7
rect 51 -1 62 7
rect -81 -108 -72 -1
rect -40 -50 75 -42
rect 88 -50 101 -42
rect -40 -89 -33 -50
rect -40 -97 -9 -89
rect 6 -97 16 -89
rect -81 -116 -9 -108
rect 6 -116 16 -108
rect -121 -133 -9 -125
rect 6 -133 17 -125
<< metal1 >>
rect -14 77 130 89
rect -6 63 1 77
rect -5 -7 1 32
rect 41 16 48 77
rect -5 -13 38 -7
rect -5 -57 1 -13
rect 78 -34 85 77
rect -5 -63 75 -57
rect -5 -78 1 -63
rect 41 -95 49 -63
rect 123 -65 130 77
rect 123 -70 156 -65
rect 41 -100 149 -95
rect 193 -99 219 -96
rect -5 -157 2 -144
rect 148 -157 156 -122
rect -9 -166 156 -157
use not  not_0
timestamp 1698771081
transform 1 0 156 0 1 -100
box -7 -28 41 38
<< labels >>
rlabel polysilicon -118 -73 -118 -73 3 a
rlabel polysilicon -77 -85 -76 -83 1 b
rlabel polysilicon -38 -83 -38 -83 1 c
rlabel metal1 91 82 92 83 1 vdd
rlabel metal1 99 -163 100 -162 1 gnd
rlabel metal1 210 -98 211 -97 1 y
<< end >>
