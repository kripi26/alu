* SPICE3 file created from decoder.ext - technology: scmos
.include TSMC_180nm.txt
.param SUPPLY = 1.8
.param LAMBDA = 0.09u
.param width_P = 8*LAMBDA
.param width_N = 4*LAMBDA
.global gnd vdd
.option scale=0.09u

Vdd vdd gnd 1.8
va0 a0 gnd pulse 0 1.8 0ns 100ps 100ps 20ns 40ns
va1 a1 gnd pulse 0 1.8 0ns 100ps 100ps 40ns 60ns


M1000 and_2/a a0 vdd not_0/vdd CMOSP w=8 l=4
+  ad=101 pd=42 as=902 ps=452
M1001 and_2/a a0 gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=866 ps=376
M1002 and_1/b a1 vdd not_1/vdd CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1003 and_1/b a1 gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1004 d0 and_0/a_n26_14# vdd and_0/vdd CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1005 vdd and_1/b and_0/a_n26_14# and_0/vdd CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1006 d0 and_0/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1007 and_0/a_n26_14# and_2/a vdd and_0/vdd CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1008 and_0/a_n26_n23# and_2/a gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1009 and_0/a_n26_14# and_1/b and_0/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1010 d1 and_1/a_n26_14# vdd and_1/vdd CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1011 vdd and_1/b and_1/a_n26_14# and_1/vdd CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1012 d1 and_1/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1013 and_1/a_n26_14# a0 vdd and_1/vdd CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1014 and_1/a_n26_n23# a0 gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1015 and_1/a_n26_14# and_1/b and_1/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1016 d2 and_2/a_n26_14# vdd and_2/vdd CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1017 vdd a1 and_2/a_n26_14# and_2/vdd CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1018 d2 and_2/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1019 and_2/a_n26_14# and_2/a vdd and_2/vdd CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1020 and_2/a_n26_n23# and_2/a gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1021 and_2/a_n26_14# a1 and_2/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1022 d3 and_3/a_n26_14# vdd and_3/vdd CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1023 vdd a1 and_3/a_n26_14# and_3/vdd CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1024 d3 and_3/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1025 and_3/a_n26_14# a0 vdd and_3/vdd CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1026 and_3/a_n26_n23# a0 gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1027 and_3/a_n26_14# a1 and_3/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
C0 and_2/vdd vdd 0.03fF
C1 vdd and_2/vdd 0.07fF
C2 a1 and_2/vdd 0.09fF
C3 d1 gnd 0.13fF
C4 vdd not_1/vdd 0.18fF
C5 a1 not_1/vdd 0.09fF
C6 and_2/a vdd 0.04fF
C7 a1 and_2/a 0.24fF
C8 d1 and_1/vdd 0.03fF
C9 and_3/a_n26_14# and_3/vdd 0.02fF
C10 a0 not_0/vdd 0.09fF
C11 and_1/b not_1/vdd 0.03fF
C12 and_2/a and_1/b 0.34fF
C13 vdd and_1/vdd 0.07fF
C14 and_0/a_n26_14# and_1/b 0.33fF
C15 gnd d2 0.14fF
C16 and_2/vdd and_2/a_n26_14# 0.09fF
C17 and_1/b and_1/vdd 0.09fF
C18 a0 and_3/vdd 0.09fF
C19 and_2/a_n26_14# and_2/vdd 0.02fF
C20 and_0/vdd and_0/a_n26_14# 0.09fF
C21 and_1/b vdd 0.04fF
C22 gnd and_2/a 0.18fF
C23 and_3/vdd vdd 0.03fF
C24 and_0/vdd vdd 0.03fF
C25 a0 and_2/a 0.12fF
C26 and_1/a_n26_14# and_1/vdd 0.02fF
C27 a1 and_3/a_n26_14# 0.31fF
C28 gnd vdd 0.80fF
C29 a1 gnd 0.34fF
C30 a1 and_2/a_n26_14# 0.31fF
C31 and_1/vdd vdd 0.03fF
C32 gnd and_1/b 0.19fF
C33 a0 and_1/vdd 0.09fF
C34 and_2/a not_0/vdd 0.03fF
C35 and_1/a_n26_14# and_1/b 0.29fF
C36 a0 vdd 0.11fF
C37 and_3/vdd and_3/a_n26_14# 0.09fF
C38 a0 a1 1.16fF
C39 and_3/vdd d3 0.03fF
C40 a0 and_1/b 0.19fF
C41 and_2/vdd d2 0.03fF
C42 and_2/a and_0/vdd 0.09fF
C43 vdd not_0/vdd 0.18fF
C44 and_0/a_n26_14# and_0/vdd 0.02fF
C45 gnd d3 0.13fF
C46 and_0/vdd d0 0.03fF
C47 and_1/a_n26_14# and_1/vdd 0.09fF
C48 gnd d0 0.01fF
C49 and_2/a and_2/vdd 0.09fF
C50 and_0/vdd vdd 0.07fF
C51 vdd and_3/vdd 0.07fF
C52 a0 gnd 0.14fF
C53 a1 and_3/vdd 0.09fF
C54 and_1/b and_0/vdd 0.09fF
C55 gnd Gnd 2.82fF
C56 d3 Gnd 0.23fF
C57 and_3/a_n26_14# Gnd 0.05fF
C58 a1 Gnd 1.05fF
C59 a0 Gnd 1.54fF
C60 vdd Gnd 4.38fF
C61 and_3/vdd Gnd 0.82fF
C62 and_3/vdd Gnd 0.82fF
C63 d2 Gnd 0.24fF
C64 and_2/a_n26_14# Gnd 0.05fF
C65 and_2/vdd Gnd 0.82fF
C66 and_2/vdd Gnd 0.82fF
C67 d1 Gnd 0.22fF
C68 and_1/a_n26_14# Gnd 0.05fF
C69 and_1/vdd Gnd 0.82fF
C70 and_1/vdd Gnd 0.82fF
C71 d0 Gnd 0.27fF
C72 and_0/a_n26_14# Gnd 0.05fF
C73 and_0/vdd Gnd 0.82fF
C74 and_0/vdd Gnd 0.82fF
C75 not_1/vdd Gnd 0.90fF
C76 not_0/vdd Gnd 0.90fF

.tran 0.1n 500n

* .measure tran trise
* + TRIG v(a) VAL = 0.9 RISE = 1
* + TARG v(out) VAL = 0.9 FALL = 1

* .measure tran tfall
* + TRIG v(a) VAL = 0.9 FALL = 1
* + TARG v(out) VAL = 0.9 RISE = 1

* .measure tran tpd param = '(trise + tfall)/2' goal = 0

.control
run
plot  v(a0) v(a1)+2 v(d0)+4 v(d1)+6 v(d2)+8 v(d3)+10
.endc

.end


