* SPICE3 file created from 4input_AND.ext - technology: scmos
.include TSMC_180nm.txt
.param SUPPLY = 1.8
.param LAMBDA = 0.09u
.param width_P = 8*LAMBDA
.param width_N = 4*LAMBDA
.global gnd vdd

Vdd vdd gnd 1.8
va a gnd pulse 0 1.8 0ns 100ps 100ps 20ns 40ns
vb b gnd pulse 0 1.8 0ns 100ps 100ps 60ns 80ns
vc c gnd pulse 0 1.8 0ns 100ps 100ps 80ns 100ns
vd d gnd pulse 0 1.8 0ns 100ps 100ps 100ns 120ns
.option scale=0.09u

M1000 y not_0/in vdd not_0/vdd CMOSP w=8 l=4
+  ad=101 pd=42 as=701 ps=238
M1001 y not_0/in gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=295 ps=98
M1002 vdd d not_0/in vdd CMOSP w=12 l=7
+  ad=0 pd=0 as=648 ps=204
M1003 not_0/in a a_n40_n132# Gnd CMOSN w=12 l=7
+  ad=120 pd=44 as=96 ps=40
M1004 a_n40_n147# c a_n40_n162# Gnd CMOSN w=12 l=7
+  ad=96 pd=40 as=96 ps=40
M1005 vdd a not_0/in vdd CMOSP w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1006 a_n40_n132# b a_n40_n147# Gnd CMOSN w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1007 a_n40_n162# d gnd Gnd CMOSN w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1008 vdd c not_0/in vdd CMOSP w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1009 vdd b not_0/in vdd CMOSP w=12 l=7
+  ad=0 pd=0 as=0 ps=0
C0 c Gnd 4.17fF
C1 d Gnd 4.88fF


.tran 0.1n 500n

* .measure tran trise
* + TRIG v(b) VAL = 0.9 RISE = 1
* + TARG v(not_0/out) VAL = 0.9 FALL = 1

* .measure tran tfall
* + TRIG v(b) VAL = 0.9 FALL = 1
* + TARG v(not_0/out) VAL = 0.9 RISE = 1

* .measure tran tpd param = '(trise + tfall)/2' goal = 0

.control
run
plot  v(a) v(b)+2 v(c)+4 v(d)+6 v(y)+8
.endc

.end



