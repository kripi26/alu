.include TSMC_180nm.txt
.include "XOR.sub"
.include "4bitadder.sub"

.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd node_x gnd 'SUPPLY'

V_in_a node_a gnd PULSE(0 1.8 0ns 100ps 100ps 180ns 200ns)
V_in_a0 node_a0 gnd PULSE(0 1.8 0ns 100ps 100ps 50ns 100ns)
V_in_a1 node_a1 gnd PULSE(0 1.8 0ns 100ps 100ps 60ns 120ns)
V_in_a2 node_a2 gnd PULSE(0 1.8 0ns 100ps 100ps 70ns 140ns)
V_in_a3 node_a3 gnd PULSE(0 1.8 0ns 100ps 100ps 80ns 160ns)
V_in_b0 node_b0 gnd PULSE(0 1.8 0ns 100ps 100ps 100ns 120ns)
V_in_b1 node_b1 gnd PULSE(0 1.8 0ns 100ps 100ps 120ns 140ns)
V_in_b2 node_b2 gnd PULSE(0 1.8 0ns 100ps 100ps 140ns 160ns)
V_in_b3 node_b3 gnd PULSE(0 1.8 0ns 100ps 100ps 160ns 180ns)

* X6 node_b0 node_a node_b0_final node_x gnd XOR
* X7 node_b1 node_a node_b1_final node_x gnd XOR
* X8 node_b2 node_a node_b2_final node_x gnd XOR
* X9 node_b3 node_a node_b3_final node_x gnd XOR

* X10 node_a0 node_b0_final node_a node_C1_add node_S0_add node_x gnd full_adder
* X11 node_a1 node_b1_final node_a node_C2_add node_S1_add node_x gnd full_adder
* X12 node_a2 node_b2_final node_a node_C3_add node_S2_add node_x gnd full_adder
* X13 node_a3 node_b3_final node_a node_C4_add node_S3_add node_x gnd full_adder

X1 node_a0 node_a1 node_a2 node_a3 node_b0 node_b1 node_b2 node_b3 gnd 5 1 2 3 4 node_x gnd 4bitadder

C1 node_C4_add gnd 100f
C2 node_S3_add gnd 100f
C3 node_S2_add gnd 100f
C4 node_S1_add gnd 100f
C5 node_S0_add gnd 100f


.tran 1n 400n


.control
run
set color0 = rgb:f/f/e
set color1 = white
plot  v(node_a) v(node_a0)+2 v(node_a1)+4 v(node_a2)+6 v(node_a3)+8
plot  v(node_b0) v(node_b1)+2 v(node_b2)+4 v(node_b3)+6
* plot  v(node_b0_final) v(node_b1_final)+2 v(node_b2_final)+4 v(node_b3_final)+6
* plot v(node_C1_add) v(node_C2_add)+2 v(node_C3_add)+4 v(node_C4_add)+6
plot v(1) v(2)+2 v(3)+4 v(4)+6 v(5)+8
* hardcopy image.ps v(node_a) v(node_b)+2 v(node_out)+4
.end
.endc

