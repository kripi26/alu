.include TSMC_180nm.txt
.include AND_block.sub

.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd node_x gnd 'SUPPLY'

V_in_a0 node_a0 gnd DC 0
V_in_a1 node_a1 gnd DC 0
V_in_a2 node_a2 gnd DC 0
V_in_a3 node_a3 gnd DC 1
V_in_b0 node_b0 gnd DC 1
V_in_b1 node_b1 gnd DC 1
V_in_b2 node_b2 gnd DC 1
V_in_b3 node_b3 gnd DC 0


X1 node_a0 node_a1 node_a2 node_a3 node_b0 node_b1 node_b2 node_b3 node_out0 node_out1 node_out2 node_out3 node_x gnd AND_block

.tran 1n 800n

C1 node_out0 gnd 100f
C2 node_out1 gnd 100f
C3 node_out2 gnd 100f
C4 node_out3 gnd 100f


.control
run
set color0 = rgb:f/f/e
set color1 = white
plot v(node_a3) v(node_a2)+2 v(node_a1)+4 v(node_a0)+6 
plot v(node_b3) v(node_b2)+2 v(node_b1)+4 v(node_b0)+6
plot v(node_out3) v(node_out2)+2 v(node_out1)+4 v(node_out0)+6

* hardcopy image.ps v(node_a) v(node_b)+2 v(node_out)+4
.end
.endc

