.include TSMC_180nm.txt
.include enable.sub

.param SUPPLY = 1.8
.param LAMBDA = 0.18u

.param wn1 = {10*LAMBDA}
.param wn2 = {10*LAMBDA}
.param ln1 = {2*LAMBDA}
.param ln2 = {2*LAMBDA}

.param wp1 = wn1
.param wp2 = wn1
.param lp1 = {LAMBDA}
.param lp2 = {LAMBDA}

.global gnd

Vdd node_x gnd 'SUPPLY'

V_in_a0 node_a0 gnd PULSE(0 1.8 0ns 100ps 100ps 20ns 50ns)
V_in_a1 node_a1 gnd PULSE(0 1.8 0ns 100ps 100ps 50ns 80ns)
V_in_a2 node_a2 gnd PULSE(0 1.8 0ns 100ps 100ps 80ns 110ns)
V_in_a3 node_a3 gnd PULSE(0 1.8 0ns 100ps 100ps 110ns 140ns)
V_in_b0 node_b0 gnd PULSE(0 1.8 0ns 100ps 100ps 140ns 180ns)
V_in_b1 node_b1 gnd PULSE(0 1.8 0ns 100ps 100ps 180ns 220ns)
V_in_b2 node_b2 gnd PULSE(0 1.8 0ns 100ps 100ps 220ns 250ns)
V_in_b3 node_b3 gnd PULSE(0 1.8 0ns 100ps 100ps 250ns 280ns)
V_in_en node_en gnd PULSE(0 1.8 0ns 100ps 100ps 280ns 320ns)

X1 node_a0 node_a1 node_a2 node_a3 node_b0 node_b1 node_b2 node_b3 node_en node_a0_out node_a1_out node_a2_out node_a3_out node_b0_out node_b1_out node_b2_out node_b3_out node_x gnd enable


.tran 1n 800n

C1 node_a0_out gnd 100f
C2 node_a1_out gnd 100f
C3 node_a2_out gnd 100f
C4 node_a3_out gnd 100f
C5 node_b0_out gnd 100f
C6 node_b1_out gnd 100f
C7 node_b2_out gnd 100f
C8 node_b3_out gnd 100f


.control
run
set color0 = rgb:f/f/e
set color1 = white
plot v(node_a3) v(node_a2)+2 v(node_a1)+4 v(node_a0)+6 v(node_en)+8
plot v(node_b3) v(node_b2)+2 v(node_b1)+4 v(node_b0)+6
plot v(node_a3_out) v(node_a2_out)+2 v(node_a1_out)+4 v(node_a0_out)+6
plot v(node_b3_out) v(node_b2_out)+2 v(node_b1_out)+4 v(node_b0_out)+6
* hardcopy image.ps v(node_a) v(node_b)+2 v(node_out)+4
.end
.endc

