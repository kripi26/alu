magic
tech scmos
timestamp 1699973769
<< nwell >>
rect -43 8 0 27
rect 26 9 69 28
<< ntransistor >>
rect -30 -23 -26 -14
rect -17 -23 -13 -14
rect 43 -24 47 -15
<< ptransistor >>
rect -30 14 -26 21
rect -17 14 -13 21
rect 43 15 47 22
<< ndiffusion >>
rect -32 -23 -30 -14
rect -26 -23 -17 -14
rect -13 -23 -10 -14
rect 36 -24 43 -15
rect 47 -24 59 -15
<< pdiffusion >>
rect -32 14 -30 21
rect -26 14 -24 21
rect -20 14 -17 21
rect -13 14 -11 21
rect 36 15 43 22
rect 47 15 59 22
<< ndcontact >>
rect -37 -23 -32 -14
rect -10 -23 -6 -14
rect 31 -24 36 -15
rect 59 -24 63 -15
<< pdcontact >>
rect -37 14 -32 21
rect -24 14 -20 21
rect -11 14 -6 21
rect 32 15 36 22
rect 59 15 63 22
<< psubstratepcontact >>
rect -31 -38 -24 -31
rect -17 -38 -10 -31
rect 0 -38 7 -31
rect 23 -38 30 -31
rect 41 -38 48 -31
rect 59 -38 66 -31
<< nsubstratencontact >>
rect -30 30 -24 36
rect -17 30 -11 36
rect -3 30 3 36
rect 17 30 23 36
rect 33 30 39 36
rect 46 30 52 36
rect 63 30 69 36
<< polysilicon >>
rect -30 21 -26 24
rect -17 21 -13 24
rect 43 22 47 25
rect -30 -14 -26 14
rect -17 -14 -13 14
rect 43 0 47 15
rect 0 -4 47 0
rect 43 -15 47 -4
rect -30 -26 -26 -23
rect -17 -26 -13 -23
rect 43 -27 47 -24
<< polycontact >>
rect -4 -4 0 0
<< metal1 >>
rect -37 30 -30 36
rect -24 30 -17 36
rect -11 30 -3 36
rect 3 30 17 36
rect 23 30 33 36
rect 39 30 46 36
rect 52 30 63 36
rect -37 21 -32 30
rect -11 21 -6 30
rect 32 22 36 30
rect -24 0 -20 14
rect -24 -4 -4 0
rect -10 -14 -6 -4
rect 59 -15 63 15
rect -37 -31 -32 -23
rect 31 -31 36 -24
rect -37 -38 -31 -31
rect -24 -38 -17 -31
rect -10 -38 0 -31
rect 7 -38 23 -31
rect 30 -38 41 -31
rect 48 -38 59 -31
rect 66 -38 74 -31
<< labels >>
rlabel metal1 -33 32 -32 33 5 vdd
rlabel metal1 -34 -35 -33 -34 1 gnd
rlabel polysilicon -29 -4 -28 -3 1 a
rlabel polysilicon -15 2 -14 3 1 b
rlabel metal1 61 -2 62 -1 1 y
<< end >>
