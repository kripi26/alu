* SPICE3 file created from comparator.ext - technology: scmos
.include TSMC_180nm.txt
.param SUPPLY = 1.8
.param LAMBDA = 0.09u
.param width_P = 8*LAMBDA
.param width_N = 4*LAMBDA
.global gnd vdd

Vdd vdd gnd 1.8
va0 a0 gnd DC 1.8
va1 a1 gnd DC 1.8
va2 a2 gnd DC 0
va3 a3 gnd DC 0
vb0 b0 gnd DC 1.8
vb1 b1 gnd DC 0
vb2 b2 gnd DC 1.8
vb3 b3 gnd DC 0

.option scale=0.09u

M1000 b0bar b0 vdd not_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=6353 ps=2634
M1001 b0bar b0 gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=10003 ps=2710
M1002 b1bar b1 vdd not_1/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1003 b1bar b1 gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1004 agb 4input_OR_0/y vdd 4input_OR_0/NOT_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1005 agb 4input_OR_0/y gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1006 vdd t8 4input_OR_0/a_n52_24# 4input_OR_0/w_n58_n43# CMOSP w=14 l=5
+  ad=0 pd=0 as=126 ps=46
M1007 4input_OR_0/y t8 gnd Gnd CMOSN w=16 l=7
+  ad=704 pd=216 as=0 ps=0
M1008 4input_OR_0/a_n52_4# t6 4input_OR_0/a_n52_n15# 4input_OR_0/w_n58_n43# CMOSP w=14 l=5
+  ad=210 pd=58 as=196 ps=56
M1009 4input_OR_0/y t5 gnd Gnd CMOSN w=16 l=7
+  ad=0 pd=0 as=0 ps=0
M1010 4input_OR_0/y t7 gnd Gnd CMOSN w=16 l=7
+  ad=0 pd=0 as=0 ps=0
M1011 4input_OR_0/a_n52_24# t7 4input_OR_0/a_n52_4# 4input_OR_0/w_n58_n43# CMOSP w=14 l=5
+  ad=0 pd=0 as=0 ps=0
M1012 4input_OR_0/a_n52_n15# t5 4input_OR_0/y 4input_OR_0/w_n58_n43# CMOSP w=14 l=5
+  ad=0 pd=0 as=238 ps=62
M1013 4input_OR_0/y t6 gnd Gnd CMOSN w=16 l=7
+  ad=0 pd=0 as=0 ps=0
M1014 b2bar b2 vdd not_2/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1015 b2bar b2 gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1016 a3xnorb3 xnor_0/not_0/in vdd xnor_0/not_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1017 a3xnorb3 xnor_0/not_0/in gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1018 xnor_0/not_0/in b3 xnor_0/XOR_0/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1019 xnor_0/XOR_0/bbar b3 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1020 xnor_0/not_0/in xnor_0/XOR_0/bbar xnor_0/XOR_0/abar xnor_0/XOR_0/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1021 vdd b3 xnor_0/XOR_0/bbar xnor_0/XOR_0/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1022 xnor_0/not_0/in b3 a3 xnor_0/XOR_0/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=72 ps=34
M1023 xnor_0/XOR_0/abar a3 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1024 vdd a3 xnor_0/XOR_0/abar xnor_0/XOR_0/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1025 xnor_0/not_0/in xnor_0/XOR_0/bbar a3 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=165 ps=52
M1026 b3bar b3 vdd not_3/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1027 b3bar b3 gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1028 a2xnorb2 xnor_1/not_0/in vdd xnor_1/not_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1029 a2xnorb2 xnor_1/not_0/in gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1030 xnor_1/not_0/in b2 xnor_1/XOR_0/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1031 xnor_1/XOR_0/bbar b2 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1032 xnor_1/not_0/in xnor_1/XOR_0/bbar xnor_1/XOR_0/abar xnor_1/XOR_0/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1033 vdd b2 xnor_1/XOR_0/bbar xnor_1/XOR_0/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1034 xnor_1/not_0/in b2 a2 xnor_1/XOR_0/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=72 ps=34
M1035 xnor_1/XOR_0/abar a2 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1036 vdd a2 xnor_1/XOR_0/abar xnor_1/XOR_0/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1037 xnor_1/not_0/in xnor_1/XOR_0/bbar a2 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=165 ps=52
M1038 a0bar a0 vdd not_4/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1039 a0bar a0 gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1040 bga 4input_OR_1/y vdd 4input_OR_1/NOT_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1041 bga 4input_OR_1/y gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1042 vdd t4 4input_OR_1/a_n52_24# 4input_OR_1/w_n58_n43# CMOSP w=14 l=5
+  ad=0 pd=0 as=126 ps=46
M1043 4input_OR_1/y t4 gnd Gnd CMOSN w=16 l=7
+  ad=704 pd=216 as=0 ps=0
M1044 4input_OR_1/a_n52_4# t2 4input_OR_1/a_n52_n15# 4input_OR_1/w_n58_n43# CMOSP w=14 l=5
+  ad=210 pd=58 as=196 ps=56
M1045 4input_OR_1/y t1 gnd Gnd CMOSN w=16 l=7
+  ad=0 pd=0 as=0 ps=0
M1046 4input_OR_1/y t3 gnd Gnd CMOSN w=16 l=7
+  ad=0 pd=0 as=0 ps=0
M1047 4input_OR_1/a_n52_24# t3 4input_OR_1/a_n52_4# 4input_OR_1/w_n58_n43# CMOSP w=14 l=5
+  ad=0 pd=0 as=0 ps=0
M1048 4input_OR_1/a_n52_n15# t1 4input_OR_1/y 4input_OR_1/w_n58_n43# CMOSP w=14 l=5
+  ad=0 pd=0 as=238 ps=62
M1049 4input_OR_1/y t2 gnd Gnd CMOSN w=16 l=7
+  ad=0 pd=0 as=0 ps=0
M1050 a1xnorb1 xnor_2/not_0/in vdd xnor_2/not_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1051 a1xnorb1 xnor_2/not_0/in gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1052 xnor_2/not_0/in b1 xnor_2/XOR_0/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1053 xnor_2/XOR_0/bbar b1 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1054 xnor_2/not_0/in xnor_2/XOR_0/bbar xnor_2/XOR_0/abar xnor_2/XOR_0/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1055 vdd b1 xnor_2/XOR_0/bbar xnor_2/XOR_0/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1056 xnor_2/not_0/in b1 a1 xnor_2/XOR_0/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=72 ps=34
M1057 xnor_2/XOR_0/abar a1 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1058 vdd a1 xnor_2/XOR_0/abar xnor_2/XOR_0/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1059 xnor_2/not_0/in xnor_2/XOR_0/bbar a1 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=165 ps=52
M1060 a0xnorb0 xnor_3/not_0/in vdd xnor_3/not_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1061 a0xnorb0 xnor_3/not_0/in gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1062 xnor_3/not_0/in b0 xnor_3/XOR_0/abar Gnd CMOSN w=11 l=6
+  ad=330 pd=104 as=407 ps=118
M1063 xnor_3/XOR_0/bbar b0 gnd Gnd CMOSN w=22 l=4
+  ad=242 pd=66 as=0 ps=0
M1064 xnor_3/not_0/in xnor_3/XOR_0/bbar xnor_3/XOR_0/abar xnor_3/XOR_0/w_62_n20# CMOSP w=12 l=6
+  ad=180 pd=76 as=218 ps=84
M1065 vdd b0 xnor_3/XOR_0/bbar xnor_3/XOR_0/w_16_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=110 ps=42
M1066 xnor_3/not_0/in b0 a0 xnor_3/XOR_0/w_62_37# CMOSP w=8 l=6
+  ad=0 pd=0 as=72 ps=34
M1067 xnor_3/XOR_0/abar a0 gnd Gnd CMOSN w=22 l=4
+  ad=0 pd=0 as=0 ps=0
M1068 vdd a0 xnor_3/XOR_0/abar xnor_3/XOR_0/w_n34_n1# CMOSP w=10 l=4
+  ad=0 pd=0 as=0 ps=0
M1069 xnor_3/not_0/in xnor_3/XOR_0/bbar a0 Gnd CMOSN w=11 l=6
+  ad=0 pd=0 as=165 ps=52
M1070 a1bar a1 vdd not_5/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1071 a1bar a1 gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1072 a2bar a2 vdd not_6/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1073 a2bar a2 gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1074 a3bar a3 vdd not_7/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1075 a3bar a3 gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1076 t8 5input_AND_0/not_0/in vdd 5input_AND_0/not_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1077 t8 5input_AND_0/not_0/in gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1078 vdd a0 5input_AND_0/not_0/in 5input_AND_0/w_n37_15# CMOSP w=14 l=8
+  ad=0 pd=0 as=405 ps=198
M1079 vdd a3xnorb3 5input_AND_0/not_0/in 5input_AND_0/w_31_n55# CMOSP w=15 l=8
+  ad=0 pd=0 as=0 ps=0
M1080 5input_AND_0/a_n33_n203# b0bar 5input_AND_0/a_n33_n226# Gnd CMOSN w=36 l=12
+  ad=468 pd=98 as=396 ps=94
M1081 5input_AND_0/not_0/in a1xnorb1 5input_AND_0/a_n33_n154# Gnd CMOSN w=36 l=12
+  ad=540 pd=102 as=432 ps=96
M1082 vdd a1xnorb1 5input_AND_0/not_0/in 5input_AND_0/w_106_n113# CMOSP w=13 l=8
+  ad=0 pd=0 as=0 ps=0
M1083 5input_AND_0/a_n33_n154# a2xnorb2 5input_AND_0/a_n33_n178# Gnd CMOSN w=36 l=12
+  ad=0 pd=0 as=432 ps=96
M1084 5input_AND_0/a_n33_n178# a3xnorb3 5input_AND_0/a_n33_n203# Gnd CMOSN w=36 l=12
+  ad=0 pd=0 as=0 ps=0
M1085 5input_AND_0/a_n33_n226# a0 gnd Gnd CMOSN w=36 l=12
+  ad=0 pd=0 as=0 ps=0
M1086 vdd b0bar 5input_AND_0/not_0/in 5input_AND_0/w_n4_n20# CMOSP w=13 l=8
+  ad=0 pd=0 as=0 ps=0
M1087 vdd a2xnorb2 5input_AND_0/not_0/in 5input_AND_0/w_68_n82# CMOSP w=14 l=8
+  ad=0 pd=0 as=0 ps=0
M1088 t4 5input_AND_1/not_0/in vdd 5input_AND_1/not_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1089 t4 5input_AND_1/not_0/in gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1090 vdd a0bar 5input_AND_1/not_0/in 5input_AND_1/w_n37_15# CMOSP w=14 l=8
+  ad=0 pd=0 as=405 ps=198
M1091 vdd a1xnorb1 5input_AND_1/not_0/in 5input_AND_1/w_31_n55# CMOSP w=15 l=8
+  ad=0 pd=0 as=0 ps=0
M1092 5input_AND_1/a_n33_n203# b0 5input_AND_1/a_n33_n226# Gnd CMOSN w=36 l=12
+  ad=468 pd=98 as=396 ps=94
M1093 5input_AND_1/not_0/in a3xnorb3 5input_AND_1/a_n33_n154# Gnd CMOSN w=36 l=12
+  ad=540 pd=102 as=432 ps=96
M1094 vdd a3xnorb3 5input_AND_1/not_0/in 5input_AND_1/w_106_n113# CMOSP w=13 l=8
+  ad=0 pd=0 as=0 ps=0
M1095 5input_AND_1/a_n33_n154# a2xnorb2 5input_AND_1/a_n33_n178# Gnd CMOSN w=36 l=12
+  ad=0 pd=0 as=432 ps=96
M1096 5input_AND_1/a_n33_n178# a1xnorb1 5input_AND_1/a_n33_n203# Gnd CMOSN w=36 l=12
+  ad=0 pd=0 as=0 ps=0
M1097 5input_AND_1/a_n33_n226# a0bar gnd Gnd CMOSN w=36 l=12
+  ad=0 pd=0 as=0 ps=0
M1098 vdd b0 5input_AND_1/not_0/in 5input_AND_1/w_n4_n20# CMOSP w=13 l=8
+  ad=0 pd=0 as=0 ps=0
M1099 vdd a2xnorb2 5input_AND_1/not_0/in 5input_AND_1/w_68_n82# CMOSP w=14 l=8
+  ad=0 pd=0 as=0 ps=0
M1100 t5 and_0/a_n26_14# vdd and_0/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1101 vdd b3bar and_0/a_n26_14# and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1102 t5 and_0/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1103 and_0/a_n26_14# a3 vdd and_0/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1104 and_0/a_n26_n23# a3 gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1105 and_0/a_n26_14# b3bar and_0/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1106 equal 4input_AND_0/not_0/in vdd 4input_AND_0/not_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1107 equal 4input_AND_0/not_0/in gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1108 vdd a3xnorb3 4input_AND_0/not_0/in 4input_AND_0/w_n47_52# CMOSP w=12 l=7
+  ad=0 pd=0 as=648 ps=204
M1109 4input_AND_0/not_0/in a0xnorb0 4input_AND_0/a_n40_n132# Gnd CMOSN w=12 l=7
+  ad=120 pd=44 as=96 ps=40
M1110 4input_AND_0/a_n40_n147# a2xnorb2 4input_AND_0/a_n40_n162# Gnd CMOSN w=12 l=7
+  ad=96 pd=40 as=96 ps=40
M1111 vdd a0xnorb0 4input_AND_0/not_0/in 4input_AND_0/w_68_n95# CMOSP w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1112 4input_AND_0/a_n40_n132# a1xnorb1 4input_AND_0/a_n40_n147# Gnd CMOSN w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1113 4input_AND_0/a_n40_n162# a3xnorb3 gnd Gnd CMOSN w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1114 vdd a2xnorb2 4input_AND_0/not_0/in 4input_AND_0/w_n8_2# CMOSP w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1115 vdd a1xnorb1 4input_AND_0/not_0/in 4input_AND_0/w_29_n46# CMOSP w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1116 t7 4input_AND_1/not_0/in vdd 4input_AND_1/not_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1117 t7 4input_AND_1/not_0/in gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1118 vdd a1 4input_AND_1/not_0/in 4input_AND_1/w_n47_52# CMOSP w=12 l=7
+  ad=0 pd=0 as=648 ps=204
M1119 4input_AND_1/not_0/in a2xnorb2 4input_AND_1/a_n40_n132# Gnd CMOSN w=12 l=7
+  ad=120 pd=44 as=96 ps=40
M1120 4input_AND_1/a_n40_n147# b1bar 4input_AND_1/a_n40_n162# Gnd CMOSN w=12 l=7
+  ad=96 pd=40 as=96 ps=40
M1121 vdd a2xnorb2 4input_AND_1/not_0/in 4input_AND_1/w_68_n95# CMOSP w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1122 4input_AND_1/a_n40_n132# a3xnorb3 4input_AND_1/a_n40_n147# Gnd CMOSN w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1123 4input_AND_1/a_n40_n162# a1 gnd Gnd CMOSN w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1124 vdd b1bar 4input_AND_1/not_0/in 4input_AND_1/w_n8_2# CMOSP w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1125 vdd a3xnorb3 4input_AND_1/not_0/in 4input_AND_1/w_29_n46# CMOSP w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1126 t1 and_1/a_n26_14# vdd and_1/w_26_9# CMOSP w=7 l=4
+  ad=112 pd=46 as=0 ps=0
M1127 vdd b3 and_1/a_n26_14# and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=63 ps=32
M1128 t1 and_1/a_n26_14# gnd Gnd CMOSN w=9 l=4
+  ad=144 pd=50 as=0 ps=0
M1129 and_1/a_n26_14# a3bar vdd and_1/w_n43_8# CMOSP w=7 l=4
+  ad=0 pd=0 as=0 ps=0
M1130 and_1/a_n26_n23# a3bar gnd Gnd CMOSN w=9 l=4
+  ad=81 pd=36 as=0 ps=0
M1131 and_1/a_n26_14# b3 and_1/a_n26_n23# Gnd CMOSN w=9 l=4
+  ad=63 pd=32 as=0 ps=0
M1132 t3 4input_AND_2/not_0/in vdd 4input_AND_2/not_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1133 t3 4input_AND_2/not_0/in gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1134 vdd a1bar 4input_AND_2/not_0/in 4input_AND_2/w_n47_52# CMOSP w=12 l=7
+  ad=0 pd=0 as=648 ps=204
M1135 4input_AND_2/not_0/in a3xnorb3 4input_AND_2/a_n40_n132# Gnd CMOSN w=12 l=7
+  ad=120 pd=44 as=96 ps=40
M1136 4input_AND_2/a_n40_n147# b1 4input_AND_2/a_n40_n162# Gnd CMOSN w=12 l=7
+  ad=96 pd=40 as=96 ps=40
M1137 vdd a3xnorb3 4input_AND_2/not_0/in 4input_AND_2/w_68_n95# CMOSP w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1138 4input_AND_2/a_n40_n132# a2xnorb2 4input_AND_2/a_n40_n147# Gnd CMOSN w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1139 4input_AND_2/a_n40_n162# a1bar gnd Gnd CMOSN w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1140 vdd b1 4input_AND_2/not_0/in 4input_AND_2/w_n8_2# CMOSP w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1141 vdd a2xnorb2 4input_AND_2/not_0/in 4input_AND_2/w_29_n46# CMOSP w=12 l=7
+  ad=0 pd=0 as=0 ps=0
M1142 t6 3input_AND_0/not_0/in vdd 3input_AND_0/not_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1143 t6 3input_AND_0/not_0/in gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1144 3input_AND_0/a_n9_n125# b2bar gnd Gnd CMOSN w=15 l=8
+  ad=135 pd=48 as=0 ps=0
M1145 3input_AND_0/not_0/in a3xnorb3 3input_AND_0/a_n9_n108# Gnd CMOSN w=15 l=8
+  ad=165 pd=52 as=165 ps=52
M1146 vdd a3xnorb3 3input_AND_0/not_0/in 3input_AND_0/w_69_n71# CMOSP w=13 l=8
+  ad=0 pd=0 as=546 ps=162
M1147 vdd a2 3input_AND_0/not_0/in 3input_AND_0/w_32_n21# CMOSP w=13 l=8
+  ad=0 pd=0 as=0 ps=0
M1148 vdd b2bar 3input_AND_0/not_0/in 3input_AND_0/w_n14_24# CMOSP w=13 l=8
+  ad=0 pd=0 as=0 ps=0
M1149 3input_AND_0/a_n9_n108# a2 3input_AND_0/a_n9_n125# Gnd CMOSN w=15 l=8
+  ad=0 pd=0 as=0 ps=0
M1150 t2 3input_AND_1/not_0/in vdd 3input_AND_1/not_0/w_n2_10# CMOSP w=8 l=4
+  ad=101 pd=42 as=0 ps=0
M1151 t2 3input_AND_1/not_0/in gnd Gnd CMOSN w=7 l=4
+  ad=84 pd=38 as=0 ps=0
M1152 3input_AND_1/a_n9_n125# a2bar gnd Gnd CMOSN w=15 l=8
+  ad=135 pd=48 as=0 ps=0
M1153 3input_AND_1/not_0/in a3xnorb3 3input_AND_1/a_n9_n108# Gnd CMOSN w=15 l=8
+  ad=165 pd=52 as=165 ps=52
M1154 vdd a3xnorb3 3input_AND_1/not_0/in 3input_AND_1/w_69_n71# CMOSP w=13 l=8
+  ad=0 pd=0 as=546 ps=162
M1155 vdd b2 3input_AND_1/not_0/in 3input_AND_1/w_32_n21# CMOSP w=13 l=8
+  ad=0 pd=0 as=0 ps=0
M1156 vdd a2bar 3input_AND_1/not_0/in 3input_AND_1/w_n14_24# CMOSP w=13 l=8
+  ad=0 pd=0 as=0 ps=0
M1157 3input_AND_1/a_n9_n108# b2 3input_AND_1/a_n9_n125# Gnd CMOSN w=15 l=8
+  ad=0 pd=0 as=0 ps=0
C0 a1 xnor_2/XOR_0/w_n34_n1# 0.11fF
C1 a2xnorb2 4input_AND_2/not_0/in 0.18fF
C2 a0 5input_AND_0/w_n37_15# 0.17fF
C3 a2xnorb2 4input_AND_0/not_0/in 0.18fF
C4 4input_AND_1/w_68_n95# vdd 0.02fF
C5 and_0/w_n43_8# and_0/a_n26_14# 0.02fF
C6 5input_AND_0/not_0/in a2xnorb2 0.23fF
C7 b3 xnor_0/XOR_0/w_16_n1# 0.11fF
C8 4input_AND_2/not_0/in gnd 0.24fF
C9 4input_AND_1/w_n47_52# 4input_AND_1/not_0/in 0.02fF
C10 4input_AND_0/not_0/in gnd 0.03fF
C11 vdd t6 0.04fF
C12 b3bar and_0/a_n26_14# 0.10fF
C13 t6 4input_OR_0/y 0.18fF
C14 5input_AND_0/not_0/in gnd 0.10fF
C15 xnor_3/not_0/in xnor_3/XOR_0/w_62_37# 0.02fF
C16 vdd a3 0.64fF
C17 4input_AND_1/w_n47_52# vdd 0.02fF
C18 and_1/a_n26_14# and_1/w_n43_8# 0.02fF
C19 4input_AND_1/w_29_n46# a3xnorb3 0.16fF
C20 5input_AND_1/w_31_n55# vdd 0.06fF
C21 b2 a3 0.17fF
C22 b1 xnor_2/XOR_0/w_16_n1# 0.11fF
C23 a1bar vdd 0.22fF
C24 5input_AND_1/w_n37_15# vdd 0.05fF
C25 not_2/w_n2_10# b2bar 0.03fF
C26 equal 4input_AND_0/not_0/w_n2_10# 0.03fF
C27 a3bar and_1/w_n43_8# 0.09fF
C28 t5 gnd 0.34fF
C29 a2bar vdd 0.45fF
C30 xnor_1/XOR_0/abar a2 0.13fF
C31 and_0/w_26_9# t5 0.03fF
C32 b1 a1 0.19fF
C33 5input_AND_0/not_0/w_n2_10# vdd 0.17fF
C34 not_7/w_n2_10# a3 0.09fF
C35 a3xnorb3 4input_AND_2/not_0/in 0.18fF
C36 a3xnorb3 4input_AND_0/w_n47_52# 0.16fF
C37 a2bar b2 0.27fF
C38 a1xnorb1 4input_AND_0/not_0/in 0.18fF
C39 equal vdd 0.04fF
C40 4input_OR_0/w_n58_n43# t8 0.13fF
C41 xnor_2/not_0/w_n2_10# a1xnorb1 0.03fF
C42 vdd xnor_1/XOR_0/w_n34_n1# 0.02fF
C43 5input_AND_0/not_0/in a3xnorb3 0.23fF
C44 5input_AND_0/not_0/in a1xnorb1 0.23fF
C45 4input_AND_1/w_n8_2# b1bar 0.16fF
C46 and_1/a_n26_14# gnd 0.02fF
C47 t7 t5 0.21fF
C48 vdd t4 0.04fF
C49 not_3/w_n2_10# b3bar 0.03fF
C50 vdd bga 0.04fF
C51 t1 t4 0.18fF
C52 a2xnorb2 5input_AND_1/not_0/in 0.23fF
C53 b0 a3 0.14fF
C54 t8 vdd 0.04fF
C55 5input_AND_1/w_68_n82# 5input_AND_1/not_0/in 0.02fF
C56 4input_OR_1/y t2 0.18fF
C57 a1xnorb1 4input_AND_0/w_29_n46# 0.16fF
C58 b1 4input_AND_2/w_n8_2# 0.16fF
C59 not_5/w_n2_10# a1 0.09fF
C60 5input_AND_1/not_0/in gnd 0.10fF
C61 xnor_1/XOR_0/bbar b2 0.02fF
C62 a2xnorb2 b3bar 0.12fF
C63 b0 xnor_3/XOR_0/abar 0.30fF
C64 4input_OR_1/y t3 0.18fF
C65 vdd xnor_1/XOR_0/w_16_n1# 0.02fF
C66 vdd b0bar 0.14fF
C67 a3xnorb3 4input_AND_2/w_n47_52# 0.04fF
C68 xnor_2/not_0/w_n2_10# xnor_2/not_0/in 0.09fF
C69 xnor_1/not_0/w_n2_10# xnor_1/not_0/in 0.09fF
C70 b3bar gnd 0.27fF
C71 vdd xnor_2/XOR_0/w_16_n1# 0.02fF
C72 xnor_1/XOR_0/w_16_n1# b2 0.11fF
C73 vdd 3input_AND_0/not_0/w_n2_10# 0.18fF
C74 5input_AND_0/w_n4_n20# b0bar 0.18fF
C75 xnor_0/XOR_0/w_62_37# a3 0.02fF
C76 5input_AND_0/w_31_n55# 5input_AND_0/not_0/in 0.03fF
C77 and_1/a_n26_14# b3 0.10fF
C78 vdd 4input_AND_0/w_n8_2# 0.02fF
C79 xnor_2/not_0/in xnor_2/XOR_0/w_62_n20# 0.04fF
C80 a2xnorb2 b2bar 0.11fF
C81 vdd a1 1.07fF
C82 not_2/w_n2_10# vdd 0.18fF
C83 a2xnorb2 b1 0.26fF
C84 vdd 5input_AND_0/w_106_n113# 0.04fF
C85 a1xnorb1 5input_AND_1/not_0/in 0.23fF
C86 a3xnorb3 5input_AND_1/not_0/in 0.23fF
C87 gnd b2bar 0.14fF
C88 3input_AND_1/w_n14_24# 3input_AND_1/not_0/in 0.03fF
C89 a1 b2 0.19fF
C90 not_2/w_n2_10# b2 0.09fF
C91 xnor_2/XOR_0/abar a1 0.13fF
C92 b1 gnd 0.71fF
C93 vdd 4input_OR_1/NOT_0/w_n2_10# 0.18fF
C94 5input_AND_1/not_0/in 5input_AND_1/not_0/w_n2_10# 0.09fF
C95 4input_AND_2/not_0/in 4input_AND_2/w_68_n95# 0.02fF
C96 vdd 4input_AND_0/w_68_n95# 0.02fF
C97 vdd xnor_3/XOR_0/w_n34_n1# 0.02fF
C98 a3xnorb3 b3bar 0.14fF
C99 xnor_0/not_0/in gnd 0.03fF
C100 5input_AND_0/not_0/in 5input_AND_0/w_n37_15# 0.05fF
C101 5input_AND_1/w_106_n113# 5input_AND_1/not_0/in 0.03fF
C102 3input_AND_1/not_0/w_n2_10# t2 0.03fF
C103 xnor_1/XOR_0/abar xnor_1/XOR_0/w_62_n20# 0.02fF
C104 vdd a0xnorb0 0.04fF
C105 xnor_2/XOR_0/bbar xnor_2/XOR_0/w_62_n20# 0.13fF
C106 vdd 4input_AND_2/w_n8_2# 0.02fF
C107 vdd xnor_3/not_0/w_n2_10# 0.18fF
C108 xnor_1/XOR_0/w_62_n20# xnor_1/not_0/in 0.04fF
C109 t8 t6 0.29fF
C110 a3xnorb3 b2bar 0.38fF
C111 vdd not_0/w_n2_10# 0.18fF
C112 5input_AND_0/w_68_n82# a2xnorb2 0.16fF
C113 not_3/w_n2_10# vdd 0.18fF
C114 a1xnorb1 b1 0.37fF
C115 a3xnorb3 b1 0.36fF
C116 vdd and_1/w_n43_8# 0.07fF
C117 b0 a1 0.19fF
C118 vdd 4input_OR_1/w_n58_n43# 0.03fF
C119 a2 b3bar 0.21fF
C120 b3 b1 0.20fF
C121 4input_AND_1/not_0/in a2xnorb2 0.18fF
C122 t6 3input_AND_0/not_0/w_n2_10# 0.03fF
C123 t1 4input_OR_1/w_n58_n43# 0.13fF
C124 b3 xnor_0/not_0/in 0.13fF
C125 a2 not_6/w_n2_10# 0.09fF
C126 t3 t2 0.19fF
C127 xnor_2/XOR_0/w_62_37# a1 0.02fF
C128 4input_AND_1/not_0/in gnd 0.21fF
C129 a2xnorb2 vdd 2.46fF
C130 5input_AND_0/not_0/w_n2_10# t8 0.03fF
C131 t7 4input_OR_0/w_n58_n43# 0.13fF
C132 5input_AND_1/w_68_n82# vdd 0.05fF
C133 a2 b2bar 0.44fF
C134 vdd gnd 3.94fF
C135 and_0/w_26_9# vdd 0.03fF
C136 4input_OR_0/y gnd 0.03fF
C137 a2 b1 0.51fF
C138 b2 gnd 0.60fF
C139 a1 a3 0.17fF
C140 4input_AND_1/w_n47_52# a1 0.16fF
C141 a0 b1 0.42fF
C142 xnor_2/not_0/in b1 0.13fF
C143 t1 gnd 0.01fF
C144 4input_AND_1/not_0/w_n2_10# 4input_AND_1/not_0/in 0.09fF
C145 xnor_2/XOR_0/abar gnd 0.14fF
C146 b0 not_0/w_n2_10# 0.09fF
C147 t7 vdd 0.04fF
C148 t7 4input_OR_0/y 0.18fF
C149 a2xnorb2 4input_AND_2/w_29_n46# 0.16fF
C150 vdd agb 0.04fF
C151 4input_AND_1/not_0/w_n2_10# vdd 0.18fF
C152 4input_AND_0/w_n47_52# 4input_AND_0/not_0/in 0.02fF
C153 4input_AND_1/not_0/in a3xnorb3 0.18fF
C154 vdd 3input_AND_0/w_32_n21# 0.03fF
C155 vdd a1xnorb1 0.87fF
C156 a3xnorb3 vdd 1.70fF
C157 xnor_3/XOR_0/abar xnor_3/XOR_0/w_n34_n1# 0.03fF
C158 not_1/w_n2_10# b1bar 0.03fF
C159 b2 3input_AND_1/not_0/in 0.19fF
C160 xnor_1/XOR_0/bbar xnor_1/XOR_0/w_16_n1# 0.03fF
C161 b0 a2xnorb2 0.69fF
C162 a1xnorb1 b2 0.10fF
C163 a3xnorb3 b2 0.19fF
C164 a0 not_4/w_n2_10# 0.09fF
C165 b3 vdd 0.47fF
C166 vdd 5input_AND_1/not_0/w_n2_10# 0.17fF
C167 xnor_3/XOR_0/w_62_n20# xnor_3/XOR_0/bbar 0.13fF
C168 b0 gnd 0.60fF
C169 a3xnorb3 3input_AND_0/w_69_n71# 0.16fF
C170 4input_AND_0/w_29_n46# 4input_AND_0/not_0/in 0.02fF
C171 b3 b2 0.18fF
C172 xnor_2/XOR_0/bbar b1 0.02fF
C173 5input_AND_1/w_106_n113# vdd 0.04fF
C174 xnor_3/XOR_0/w_16_n1# vdd 0.02fF
C175 4input_AND_1/w_68_n95# a2xnorb2 0.16fF
C176 b3 xnor_0/XOR_0/bbar 0.02fF
C177 4input_AND_2/not_0/in 4input_AND_2/w_n47_52# 0.02fF
C178 bga 4input_OR_1/NOT_0/w_n2_10# 0.03fF
C179 3input_AND_1/w_32_n21# 3input_AND_1/not_0/in 0.02fF
C180 3input_AND_0/not_0/in 3input_AND_0/w_n14_24# 0.03fF
C181 4input_AND_2/not_0/w_n2_10# t3 0.03fF
C182 vdd a2 1.34fF
C183 3input_AND_0/not_0/in 3input_AND_0/w_69_n71# 0.02fF
C184 a2xnorb2 a3 0.15fF
C185 a0 vdd 0.49fF
C186 a2 b2 0.17fF
C187 xnor_0/XOR_0/abar xnor_0/XOR_0/w_62_n20# 0.02fF
C188 4input_AND_2/not_0/in 4input_AND_2/not_0/w_n2_10# 0.09fF
C189 5input_AND_0/w_31_n55# vdd 0.06fF
C190 a0 b2 0.16fF
C191 b0 a1xnorb1 0.51fF
C192 b0 a3xnorb3 0.48fF
C193 5input_AND_1/w_n4_n20# 5input_AND_1/not_0/in 0.03fF
C194 a1bar a2xnorb2 0.26fF
C195 a3 gnd 0.43fF
C196 xnor_0/not_0/w_n2_10# a3xnorb3 0.03fF
C197 xnor_3/XOR_0/w_62_n20# xnor_3/not_0/in 0.04fF
C198 4input_AND_1/w_n8_2# 4input_AND_1/not_0/in 0.02fF
C199 t7 t6 0.27fF
C200 b0 b3 0.15fF
C201 vdd xnor_0/XOR_0/w_n34_n1# 0.02fF
C202 4input_OR_1/w_n58_n43# t4 0.13fF
C203 t1 4input_OR_1/y 0.18fF
C204 a0bar not_4/w_n2_10# 0.03fF
C205 xnor_3/XOR_0/abar gnd 0.14fF
C206 4input_AND_1/w_n8_2# vdd 0.02fF
C207 4input_OR_0/NOT_0/w_n2_10# vdd 0.18fF
C208 4input_OR_0/NOT_0/w_n2_10# 4input_OR_0/y 0.09fF
C209 xnor_3/XOR_0/w_16_n1# b0 0.11fF
C210 vdd xnor_1/not_0/w_n2_10# 0.18fF
C211 vdd 5input_AND_0/w_n37_15# 0.05fF
C212 not_0/w_n2_10# b0bar 0.03fF
C213 vdd 4input_AND_2/w_68_n95# 0.02fF
C214 xnor_0/XOR_0/abar a3 0.13fF
C215 b0 xnor_3/XOR_0/w_62_37# 0.13fF
C216 a3xnorb3 a3 0.18fF
C217 a1xnorb1 a3 0.17fF
C218 b0 a2 0.17fF
C219 b3 xnor_0/XOR_0/w_62_37# 0.13fF
C220 3input_AND_1/w_69_n71# vdd 0.03fF
C221 5input_AND_1/w_31_n55# a1xnorb1 0.21fF
C222 b0 a0 0.38fF
C223 4input_AND_1/not_0/in b1bar 0.18fF
C224 xnor_1/XOR_0/w_62_37# a2 0.02fF
C225 b3 a3 3.02fF
C226 a1bar a3xnorb3 0.36fF
C227 4input_AND_2/not_0/in b1 0.18fF
C228 vdd a0bar 0.30fF
C229 b1bar vdd 0.20fF
C230 a0xnorb0 4input_AND_0/w_68_n95# 0.16fF
C231 a2bar a3xnorb3 0.19fF
C232 xnor_2/XOR_0/w_62_37# xnor_2/not_0/in 0.02fF
C233 a2xnorb2 b0bar 0.38fF
C234 b0 xnor_3/XOR_0/bbar 0.02fF
C235 vdd 3input_AND_1/not_0/w_n2_10# 0.18fF
C236 t7 t8 0.15fF
C237 vdd xnor_0/XOR_0/w_16_n1# 0.02fF
C238 a2xnorb2 4input_AND_0/w_n8_2# 0.16fF
C239 a0xnorb0 xnor_3/not_0/w_n2_10# 0.03fF
C240 a2 a3 0.17fF
C241 a0 a3 0.10fF
C242 xnor_1/XOR_0/abar b2 0.30fF
C243 4input_AND_1/w_29_n46# 4input_AND_1/not_0/in 0.02fF
C244 a2xnorb2 a1 0.61fF
C245 5input_AND_1/not_0/w_n2_10# t4 0.03fF
C246 xnor_0/XOR_0/bbar xnor_0/XOR_0/w_16_n1# 0.03fF
C247 b2 xnor_1/not_0/in 0.13fF
C248 and_0/a_n26_14# gnd 0.00fF
C249 vdd t2 0.04fF
C250 a0 xnor_3/XOR_0/abar 0.13fF
C251 4input_AND_1/w_29_n46# vdd 0.02fF
C252 a1 gnd 0.52fF
C253 and_0/w_26_9# and_0/a_n26_14# 0.09fF
C254 and_0/w_n43_8# b3bar 0.09fF
C255 xnor_0/XOR_0/w_n34_n1# a3 0.11fF
C256 5input_AND_0/w_68_n82# 5input_AND_0/not_0/in 0.02fF
C257 b0 a0bar 0.33fF
C258 b0 xnor_3/not_0/in 0.13fF
C259 t1 t2 0.18fF
C260 a3xnorb3 b0bar 0.28fF
C261 a1xnorb1 b0bar 0.29fF
C262 vdd t3 0.04fF
C263 xnor_1/XOR_0/w_n34_n1# a2 0.11fF
C264 4input_AND_0/not_0/w_n2_10# 4input_AND_0/not_0/in 0.09fF
C265 and_1/a_n26_14# and_1/w_26_9# 0.09fF
C266 a2xnorb2 a0xnorb0 0.36fF
C267 5input_AND_1/w_n4_n20# vdd 0.05fF
C268 vdd 4input_AND_0/w_n47_52# 0.02fF
C269 t1 t3 0.18fF
C270 xnor_2/not_0/w_n2_10# vdd 0.18fF
C271 a0xnorb0 gnd 0.36fF
C272 4input_OR_0/w_n58_n43# t5 0.13fF
C273 not_1/w_n2_10# b1 0.09fF
C274 a1xnorb1 a1 0.19fF
C275 a3xnorb3 a1 0.53fF
C276 5input_AND_0/not_0/in 5input_AND_0/w_n4_n20# 0.03fF
C277 a1xnorb1 5input_AND_0/w_106_n113# 0.17fF
C278 3input_AND_0/not_0/in 3input_AND_0/not_0/w_n2_10# 0.09fF
C279 xnor_1/XOR_0/w_62_37# xnor_1/not_0/in 0.02fF
C280 b3 a1 0.18fF
C281 xnor_2/XOR_0/abar xnor_2/XOR_0/w_62_n20# 0.02fF
C282 4input_AND_2/not_0/in 4input_AND_2/w_29_n46# 0.02fF
C283 vdd 4input_AND_0/w_29_n46# 0.02fF
C284 a0 b0bar 0.25fF
C285 4input_OR_0/y t5 0.18fF
C286 5input_AND_1/w_n37_15# a0bar 0.17fF
C287 5input_AND_1/w_68_n82# a2xnorb2 0.16fF
C288 a3xnorb3 a0xnorb0 0.29fF
C289 a0xnorb0 a1xnorb1 0.40fF
C290 vdd 4input_AND_2/w_n47_52# 0.02fF
C291 5input_AND_1/w_n4_n20# b0 0.18fF
C292 a2xnorb2 gnd 1.27fF
C293 a2 a1 0.31fF
C294 a0 a1 0.13fF
C295 vdd 4input_AND_2/not_0/w_n2_10# 0.18fF
C296 a3bar vdd 0.04fF
C297 vdd xnor_2/XOR_0/w_n34_n1# 0.02fF
C298 not_3/w_n2_10# b3 0.09fF
C299 a0 xnor_3/XOR_0/w_n34_n1# 0.11fF
C300 b3 and_1/w_n43_8# 0.09fF
C301 vdd 3input_AND_1/w_n14_24# 0.03fF
C302 4input_OR_1/y 4input_OR_1/NOT_0/w_n2_10# 0.09fF
C303 and_0/w_n43_8# vdd 0.07fF
C304 xnor_1/XOR_0/abar xnor_1/XOR_0/w_n34_n1# 0.03fF
C305 xnor_2/XOR_0/abar xnor_2/XOR_0/w_n34_n1# 0.03fF
C306 xnor_2/XOR_0/bbar xnor_2/XOR_0/w_16_n1# 0.03fF
C307 not_1/w_n2_10# vdd 0.18fF
C308 a3xnorb3 a2xnorb2 7.69fF
C309 a2xnorb2 a1xnorb1 1.39fF
C310 vdd b3bar 0.04fF
C311 a3bar not_7/w_n2_10# 0.03fF
C312 gnd 3input_AND_1/not_0/in 0.21fF
C313 xnor_0/XOR_0/abar gnd 0.14fF
C314 a3xnorb3 gnd 0.82fF
C315 a1xnorb1 gnd 0.87fF
C316 vdd not_6/w_n2_10# 0.18fF
C317 4input_AND_1/not_0/w_n2_10# t7 0.03fF
C318 t4 t2 0.19fF
C319 b3 gnd 0.67fF
C320 vdd b2bar 1.10fF
C321 t6 t5 0.21fF
C322 t3 t4 0.19fF
C323 xnor_1/XOR_0/bbar xnor_1/XOR_0/w_62_n20# 0.13fF
C324 vdd b1 1.08fF
C325 4input_OR_1/y 4input_OR_1/w_n58_n43# 0.02fF
C326 b2bar 3input_AND_0/w_n14_24# 0.16fF
C327 b1bar a1 0.18fF
C328 3input_AND_0/not_0/in gnd 0.21fF
C329 5input_AND_0/not_0/in 5input_AND_0/not_0/w_n2_10# 0.09fF
C330 b0 5input_AND_1/not_0/in 0.23fF
C331 b1 b2 0.22fF
C332 a2xnorb2 a2 0.17fF
C333 a0 a2xnorb2 0.38fF
C334 a3xnorb3 3input_AND_1/not_0/in 0.19fF
C335 xnor_2/XOR_0/abar b1 0.30fF
C336 a3xnorb3 a1xnorb1 1.11fF
C337 a2 gnd 0.61fF
C338 vdd and_1/w_26_9# 0.03fF
C339 xnor_2/not_0/in gnd 0.03fF
C340 a0 gnd 0.17fF
C341 b3 xnor_0/XOR_0/abar 0.30fF
C342 b3 a1xnorb1 0.19fF
C343 a1bar 4input_AND_2/w_n47_52# 0.16fF
C344 4input_OR_1/y gnd 0.03fF
C345 3input_AND_0/not_0/in 3input_AND_0/w_32_n21# 0.02fF
C346 t1 and_1/w_26_9# 0.03fF
C347 5input_AND_1/w_106_n113# a3xnorb3 0.17fF
C348 not_5/w_n2_10# vdd 0.18fF
C349 vdd not_4/w_n2_10# 0.26fF
C350 xnor_3/not_0/in xnor_3/not_0/w_n2_10# 0.09fF
C351 3input_AND_0/not_0/in a3xnorb3 0.19fF
C352 5input_AND_0/w_68_n82# vdd 0.05fF
C353 a2 3input_AND_0/w_32_n21# 0.16fF
C354 4input_OR_0/w_n58_n43# vdd 0.03fF
C355 5input_AND_1/w_31_n55# 5input_AND_1/not_0/in 0.03fF
C356 a2xnorb2 xnor_1/not_0/w_n2_10# 0.03fF
C357 5input_AND_0/not_0/in b0bar 0.23fF
C358 4input_OR_0/w_n58_n43# 4input_OR_0/y 0.02fF
C359 b0 b1 0.41fF
C360 and_0/w_n43_8# a3 0.09fF
C361 a1xnorb1 a2 0.17fF
C362 a3xnorb3 a2 0.60fF
C363 xnor_0/not_0/in xnor_0/XOR_0/w_62_n20# 0.04fF
C364 t8 t5 0.21fF
C365 4input_AND_0/w_n8_2# 4input_AND_0/not_0/in 0.02fF
C366 a0 a3xnorb3 0.28fF
C367 a0 a1xnorb1 0.40fF
C368 a3 b3bar 3.31fF
C369 vdd 4input_AND_0/not_0/w_n2_10# 0.18fF
C370 5input_AND_1/w_n37_15# 5input_AND_1/not_0/in 0.05fF
C371 xnor_0/not_0/w_n2_10# xnor_0/not_0/in 0.09fF
C372 5input_AND_0/w_31_n55# a3xnorb3 0.21fF
C373 b3 a2 0.17fF
C374 a0 b3 0.11fF
C375 a2xnorb2 a0bar 0.41fF
C376 xnor_2/XOR_0/w_62_37# b1 0.13fF
C377 a2bar 3input_AND_1/w_n14_24# 0.16fF
C378 4input_OR_0/NOT_0/w_n2_10# agb 0.03fF
C379 b1bar a2xnorb2 0.51fF
C380 xnor_0/XOR_0/abar xnor_0/XOR_0/w_n34_n1# 0.03fF
C381 vdd b2 1.23fF
C382 5input_AND_0/not_0/in 5input_AND_0/w_106_n113# 0.03fF
C383 vdd 5input_AND_0/w_n4_n20# 0.05fF
C384 3input_AND_0/not_0/in a2 0.19fF
C385 vdd 3input_AND_0/w_n14_24# 0.03fF
C386 b1bar gnd 0.14fF
C387 xnor_3/not_0/in gnd 0.03fF
C388 vdd 3input_AND_0/w_69_n71# 0.03fF
C389 4input_AND_0/w_68_n95# 4input_AND_0/not_0/in 0.02fF
C390 xnor_0/not_0/in xnor_0/XOR_0/w_62_37# 0.02fF
C391 b1 a3 0.19fF
C392 a2bar not_6/w_n2_10# 0.03fF
C393 a0 xnor_3/XOR_0/w_62_37# 0.02fF
C394 vdd not_7/w_n2_10# 0.26fF
C395 4input_OR_1/w_n58_n43# t2 0.13fF
C396 a0 a2 0.17fF
C397 4input_AND_2/not_0/in 4input_AND_2/w_n8_2# 0.02fF
C398 a3xnorb3 4input_AND_2/w_68_n95# 0.16fF
C399 vdd 4input_AND_2/w_29_n46# 0.02fF
C400 a0xnorb0 4input_AND_0/not_0/in 0.18fF
C401 a1bar b1 0.44fF
C402 xnor_3/XOR_0/w_16_n1# xnor_3/XOR_0/bbar 0.03fF
C403 3input_AND_1/w_69_n71# 3input_AND_1/not_0/in 0.02fF
C404 3input_AND_1/w_32_n21# vdd 0.03fF
C405 xnor_1/XOR_0/abar gnd 0.14fF
C406 a3xnorb3 3input_AND_1/w_69_n71# 0.16fF
C407 4input_OR_1/w_n58_n43# t3 0.13fF
C408 3input_AND_1/w_32_n21# b2 0.16fF
C409 xnor_1/not_0/in gnd 0.03fF
C410 a1xnorb1 a0bar 0.03fF
C411 a3xnorb3 a0bar 0.29fF
C412 b0 vdd 0.73fF
C413 b1bar a3xnorb3 0.35fF
C414 xnor_0/not_0/w_n2_10# vdd 0.18fF
C415 xnor_3/XOR_0/w_62_n20# xnor_3/XOR_0/abar 0.02fF
C416 3input_AND_1/not_0/w_n2_10# 3input_AND_1/not_0/in 0.09fF
C417 b0 b2 0.16fF
C418 4input_OR_0/w_n58_n43# t6 0.13fF
C419 4input_AND_1/w_68_n95# 4input_AND_1/not_0/in 0.02fF
C420 xnor_1/XOR_0/w_62_37# b2 0.13fF
C421 not_5/w_n2_10# a1bar 0.03fF
C422 xnor_0/XOR_0/bbar xnor_0/XOR_0/w_62_n20# 0.13fF
C423 a2bar Gnd 5.34fF
C424 3input_AND_1/w_69_n71# Gnd 1.13fF
C425 3input_AND_1/w_32_n21# Gnd 1.13fF
C426 3input_AND_1/w_n14_24# Gnd 1.13fF
C427 gnd Gnd 142.74fF
C428 t2 Gnd 3.00fF
C429 3input_AND_1/not_0/in Gnd 1.59fF
C430 3input_AND_1/not_0/w_n2_10# Gnd 0.90fF
C431 b2bar Gnd 5.92fF
C432 3input_AND_0/w_69_n71# Gnd 1.13fF
C433 3input_AND_0/w_32_n21# Gnd 1.13fF
C434 3input_AND_0/w_n14_24# Gnd 1.13fF
C435 t6 Gnd 2.94fF
C436 3input_AND_0/not_0/in Gnd 1.59fF
C437 3input_AND_0/not_0/w_n2_10# Gnd 0.90fF
C438 a2xnorb2 Gnd 18.99fF
C439 4input_AND_2/w_68_n95# Gnd 1.13fF
C440 4input_AND_2/w_29_n46# Gnd 1.13fF
C441 4input_AND_2/w_n8_2# Gnd 1.13fF
C442 4input_AND_2/w_n47_52# Gnd 1.13fF
C443 t3 Gnd 4.44fF
C444 4input_AND_2/not_0/in Gnd 2.38fF
C445 4input_AND_2/not_0/w_n2_10# Gnd 0.90fF
C446 and_1/a_n26_14# Gnd 0.05fF
C447 a3bar Gnd 4.39fF
C448 and_1/w_26_9# Gnd 0.82fF
C449 and_1/w_n43_8# Gnd 0.82fF
C450 4input_AND_1/w_68_n95# Gnd 1.13fF
C451 4input_AND_1/w_29_n46# Gnd 1.13fF
C452 4input_AND_1/w_n8_2# Gnd 1.13fF
C453 4input_AND_1/w_n47_52# Gnd 1.13fF
C454 t7 Gnd 4.39fF
C455 4input_AND_1/not_0/in Gnd 2.38fF
C456 4input_AND_1/not_0/w_n2_10# Gnd 0.90fF
C457 4input_AND_0/w_68_n95# Gnd 1.13fF
C458 4input_AND_0/w_29_n46# Gnd 1.13fF
C459 4input_AND_0/w_n8_2# Gnd 1.13fF
C460 4input_AND_0/w_n47_52# Gnd 1.13fF
C461 equal Gnd 0.15fF
C462 4input_AND_0/not_0/in Gnd 2.38fF
C463 4input_AND_0/not_0/w_n2_10# Gnd 0.90fF
C464 and_0/a_n26_14# Gnd 0.05fF
C465 b3bar Gnd 0.68fF
C466 and_0/w_26_9# Gnd 0.82fF
C467 and_0/w_n43_8# Gnd 0.82fF
C468 5input_AND_1/w_106_n113# Gnd 0.81fF
C469 5input_AND_1/w_68_n82# Gnd 0.81fF
C470 5input_AND_1/w_31_n55# Gnd 1.18fF
C471 5input_AND_1/w_n4_n20# Gnd 0.89fF
C472 5input_AND_1/w_n37_15# Gnd 0.89fF
C473 t4 Gnd 2.77fF
C474 5input_AND_1/not_0/in Gnd 2.73fF
C475 5input_AND_1/not_0/w_n2_10# Gnd 0.90fF
C476 5input_AND_0/w_106_n113# Gnd 0.81fF
C477 5input_AND_0/w_68_n82# Gnd 0.81fF
C478 5input_AND_0/w_31_n55# Gnd 1.18fF
C479 5input_AND_0/w_n4_n20# Gnd 0.89fF
C480 5input_AND_0/w_n37_15# Gnd 0.89fF
C481 t8 Gnd 1.96fF
C482 5input_AND_0/not_0/in Gnd 2.73fF
C483 5input_AND_0/not_0/w_n2_10# Gnd 0.90fF
C484 not_7/w_n2_10# Gnd 0.90fF
C485 not_6/w_n2_10# Gnd 0.90fF
C486 a1bar Gnd 5.03fF
C487 not_5/w_n2_10# Gnd 0.90fF
C488 xnor_3/XOR_0/abar Gnd 0.11fF
C489 xnor_3/XOR_0/bbar Gnd 0.06fF
C490 xnor_3/not_0/in Gnd 0.39fF
C491 b0 Gnd 8.34fF
C492 a0 Gnd 31.80fF
C493 xnor_3/XOR_0/w_62_n20# Gnd 0.87fF
C494 xnor_3/XOR_0/w_16_n1# Gnd 0.75fF
C495 xnor_3/XOR_0/w_n34_n1# Gnd 0.75fF
C496 xnor_3/XOR_0/w_62_37# Gnd 0.72fF
C497 a0xnorb0 Gnd 2.96fF
C498 xnor_3/not_0/w_n2_10# Gnd 0.90fF
C499 xnor_2/XOR_0/abar Gnd 0.11fF
C500 xnor_2/XOR_0/bbar Gnd 0.06fF
C501 xnor_2/not_0/in Gnd 0.39fF
C502 b1 Gnd 54.66fF
C503 a1 Gnd 41.48fF
C504 xnor_2/XOR_0/w_62_n20# Gnd 0.87fF
C505 xnor_2/XOR_0/w_16_n1# Gnd 0.75fF
C506 xnor_2/XOR_0/w_n34_n1# Gnd 0.75fF
C507 xnor_2/XOR_0/w_62_37# Gnd 0.72fF
C508 xnor_2/not_0/w_n2_10# Gnd 0.90fF
C509 4input_OR_1/w_n58_n43# Gnd 2.55fF
C510 bga Gnd 0.12fF
C511 4input_OR_1/y Gnd 1.46fF
C512 4input_OR_1/NOT_0/w_n2_10# Gnd 0.90fF
C513 a0bar Gnd 6.16fF
C514 not_4/w_n2_10# Gnd 0.90fF
C515 xnor_1/XOR_0/abar Gnd 0.11fF
C516 xnor_1/XOR_0/bbar Gnd 0.06fF
C517 xnor_1/not_0/in Gnd 0.39fF
C518 b2 Gnd 46.25fF
C519 a2 Gnd 27.53fF
C520 xnor_1/XOR_0/w_62_n20# Gnd 0.87fF
C521 xnor_1/XOR_0/w_16_n1# Gnd 0.75fF
C522 xnor_1/XOR_0/w_n34_n1# Gnd 0.75fF
C523 xnor_1/XOR_0/w_62_37# Gnd 0.72fF
C524 xnor_1/not_0/w_n2_10# Gnd 0.90fF
C525 not_3/w_n2_10# Gnd 0.90fF
C526 xnor_0/XOR_0/abar Gnd 0.11fF
C527 xnor_0/XOR_0/bbar Gnd 0.06fF
C528 xnor_0/not_0/in Gnd 0.39fF
C529 b3 Gnd 29.34fF
C530 a3 Gnd 20.52fF
C531 xnor_0/XOR_0/w_62_n20# Gnd 0.87fF
C532 xnor_0/XOR_0/w_16_n1# Gnd 0.75fF
C533 xnor_0/XOR_0/w_n34_n1# Gnd 0.75fF
C534 xnor_0/XOR_0/w_62_37# Gnd 0.72fF
C535 xnor_0/not_0/w_n2_10# Gnd 0.90fF
C536 not_2/w_n2_10# Gnd 0.90fF
C537 4input_OR_0/w_n58_n43# Gnd 2.55fF
C538 agb Gnd 0.11fF
C539 4input_OR_0/y Gnd 1.46fF
C540 vdd Gnd 81.67fF
C541 4input_OR_0/NOT_0/w_n2_10# Gnd 0.90fF
C542 b1bar Gnd 4.66fF
C543 not_1/w_n2_10# Gnd 0.90fF
C544 b0bar Gnd 6.97fF
C545 not_0/w_n2_10# Gnd 0.90fF
.tran 0.1n 100n

.control
run
plot v(a0) v(a1)+2 v(a2)+4 v(a3)+6
plot v(b0) v(b1)+2 v(b2)+4 v(b3)+6
* plot v(t1) v(t2)+2 v(t3)+4 v(t4)+6
plot  v(equal) v(agb)+2 v(bga)+4
.endc
.end
