magic
tech scmos
timestamp 1700455425
<< nwell >>
rect -48 101 43 129
rect 58 101 113 129
<< ntransistor >>
rect -20 32 -15 48
rect 4 32 9 48
rect 83 32 89 48
<< ptransistor >>
rect -20 107 -15 123
rect 4 107 9 123
rect 83 107 89 123
<< ndiffusion >>
rect -42 42 -20 48
rect -34 32 -20 42
rect -15 38 -9 48
rect -1 38 4 48
rect -15 32 4 38
rect 9 42 37 48
rect 9 32 29 42
rect 66 41 83 48
rect 73 32 83 41
rect 89 36 99 48
rect 105 36 109 48
rect 89 32 109 36
<< pdiffusion >>
rect -33 107 -20 123
rect -15 107 4 123
rect 9 107 28 123
rect 71 107 83 123
rect 89 121 107 123
rect 89 107 99 121
rect 105 107 107 121
<< ndcontact >>
rect -42 32 -34 42
rect -9 38 -1 48
rect 29 32 37 42
rect 66 32 73 41
rect 99 36 105 48
<< pdcontact >>
rect -42 107 -33 123
rect 28 107 37 123
rect 64 107 71 123
rect 99 107 105 121
<< psubstratepcontact >>
rect -32 0 -24 7
rect -7 0 1 7
rect 18 0 26 7
<< nsubstratencontact >>
rect -30 152 -22 161
rect -7 152 1 161
rect 15 152 23 161
rect 46 152 54 161
<< polysilicon >>
rect -20 123 -15 136
rect 4 123 9 136
rect 83 123 89 140
rect -20 48 -15 107
rect 4 48 9 107
rect 83 92 89 107
rect 65 86 89 92
rect 83 48 89 86
rect -20 22 -15 32
rect 4 22 9 32
rect 83 22 89 32
<< polycontact >>
rect 59 86 65 92
<< metal1 >>
rect -42 152 -30 161
rect -22 152 -7 161
rect 1 152 15 161
rect 23 152 46 161
rect 54 152 71 161
rect -42 123 -33 152
rect 64 123 71 152
rect 28 92 37 107
rect 28 86 59 92
rect 28 79 37 86
rect -9 70 37 79
rect 99 81 105 107
rect 99 75 125 81
rect -9 48 -1 70
rect 99 48 105 75
rect -42 7 -34 32
rect 29 7 37 32
rect 66 7 73 32
rect -42 0 -32 7
rect -24 0 -7 7
rect 1 0 18 7
rect 26 0 73 7
<< labels >>
rlabel metal1 -12 155 -11 157 5 vdd
rlabel metal1 1 1 2 3 1 gnd
rlabel polysilicon -19 88 -18 90 1 a
rlabel polysilicon 5 88 6 90 1 b
rlabel metal1 115 77 116 79 1 y
<< end >>
